`ifndef SIMON_SEQ_LIST
`define SIMON_SEQ_LIST

package simon_seq_list;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import simon_agent_pkg::*;
  import simon_ref_model_pkg::*;
  import simon_env_pkg::*;

  //including simon test list

  `include "simon_basic_seq.sv"

endpackage
`endif
