/home/t/Desktop/xsim_verif_example/Adder_4_bit/src/design/half_adder.sv