module simon128s192_enc (
  input wire clk,
  input wire rst
);

endmodule
