package simon_macros;
  
  
endpackage