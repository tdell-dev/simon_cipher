  module simon128s128_enc (
    input wire clk,
    input wire rst
  );


  endmodule
