module simon96s96_enc (
  input wire clk,
  input wire rst
  );

  endmodule
