//NOTE THIS FILE IS FOR SIMULATION ONLY
`timescale 1ns / 1ps
module simon_key_bram (
  input wire clka,
  input wire ena,
  input wire wea,
  input wire [8:0] addra,
  input wire [63:0] dina,

  input wire clkb,
  input wire enb,
  input wire [8:0]  addrb,
  output logic [63:0] doutb
);

//There are 512 entries, expand it out
logic [511:0][63:0] mem_space;
logic [63:0] doutb_pipe;
logic [ 8:0] addr_store;

always_ff@(posedge clka) begin
  if ( ena & wea ) begin
    case ( addra ) 
      9'd0: begin
        mem_space[0] <= dina;
      end 
      9'd1: begin
        mem_space[1] <= dina;
      end 
      9'd2: begin
        mem_space[2] <= dina;
      end 
      9'd3: begin
        mem_space[3] <= dina;
      end 
      9'd4: begin
        mem_space[4] <= dina;
      end 
      9'd5: begin
        mem_space[5] <= dina;
      end 
      9'd6: begin
        mem_space[6] <= dina;
      end 
      9'd7: begin
        mem_space[7] <= dina;
      end 
      9'd8: begin
        mem_space[8] <= dina;
      end 
      9'd9: begin
        mem_space[9] <= dina;
      end 
      9'd10: begin
        mem_space[10] <= dina;
      end 
      9'd11: begin
        mem_space[11] <= dina;
      end 
      9'd12: begin
        mem_space[12] <= dina;
      end 
      9'd13: begin
        mem_space[13] <= dina;
      end 
      9'd14: begin
        mem_space[14] <= dina;
      end 
      9'd15: begin
        mem_space[15] <= dina;
      end 
      9'd16: begin
        mem_space[16] <= dina;
      end 
      9'd17: begin
        mem_space[17] <= dina;
      end 
      9'd18: begin
        mem_space[18] <= dina;
      end 
      9'd19: begin
        mem_space[19] <= dina;
      end 
      9'd20: begin
        mem_space[20] <= dina;
      end 
      9'd21: begin
        mem_space[21] <= dina;
      end 
      9'd22: begin
        mem_space[22] <= dina;
      end 
      9'd23: begin
        mem_space[23] <= dina;
      end 
      9'd24: begin
        mem_space[24] <= dina;
      end 
      9'd25: begin
        mem_space[25] <= dina;
      end 
      9'd26: begin
        mem_space[26] <= dina;
      end 
      9'd27: begin
        mem_space[27] <= dina;
      end 
      9'd28: begin
        mem_space[28] <= dina;
      end 
      9'd29: begin
        mem_space[29] <= dina;
      end 
      9'd30: begin
        mem_space[30] <= dina;
      end 
      9'd31: begin
        mem_space[31] <= dina;
      end 
      9'd32: begin
        mem_space[32] <= dina;
      end 
      9'd33: begin
        mem_space[33] <= dina;
      end 
      9'd34: begin
        mem_space[34] <= dina;
      end 
      9'd35: begin
        mem_space[35] <= dina;
      end 
      9'd36: begin
        mem_space[36] <= dina;
      end 
      9'd37: begin
        mem_space[37] <= dina;
      end 
      9'd38: begin
        mem_space[38] <= dina;
      end 
      9'd39: begin
        mem_space[39] <= dina;
      end 
      9'd40: begin
        mem_space[40] <= dina;
      end 
      9'd41: begin
        mem_space[41] <= dina;
      end 
      9'd42: begin
        mem_space[42] <= dina;
      end 
      9'd43: begin
        mem_space[43] <= dina;
      end 
      9'd44: begin
        mem_space[44] <= dina;
      end 
      9'd45: begin
        mem_space[45] <= dina;
      end 
      9'd46: begin
        mem_space[46] <= dina;
      end 
      9'd47: begin
        mem_space[47] <= dina;
      end 
      9'd48: begin
        mem_space[48] <= dina;
      end 
      9'd49: begin
        mem_space[49] <= dina;
      end 
      9'd50: begin
        mem_space[50] <= dina;
      end 
      9'd51: begin
        mem_space[51] <= dina;
      end 
      9'd52: begin
        mem_space[52] <= dina;
      end 
      9'd53: begin
        mem_space[53] <= dina;
      end 
      9'd54: begin
        mem_space[54] <= dina;
      end 
      9'd55: begin
        mem_space[55] <= dina;
      end 
      9'd56: begin
        mem_space[56] <= dina;
      end 
      9'd57: begin
        mem_space[57] <= dina;
      end 
      9'd58: begin
        mem_space[58] <= dina;
      end 
      9'd59: begin
        mem_space[59] <= dina;
      end 
      9'd60: begin
        mem_space[60] <= dina;
      end 
      9'd61: begin
        mem_space[61] <= dina;
      end 
      9'd62: begin
        mem_space[62] <= dina;
      end 
      9'd63: begin
        mem_space[63] <= dina;
      end 
      9'd64: begin
        mem_space[64] <= dina;
      end 
      9'd65: begin
        mem_space[65] <= dina;
      end 
      9'd66: begin
        mem_space[66] <= dina;
      end 
      9'd67: begin
        mem_space[67] <= dina;
      end 
      9'd68: begin
        mem_space[68] <= dina;
      end 
      9'd69: begin
        mem_space[69] <= dina;
      end 
      9'd70: begin
        mem_space[70] <= dina;
      end 
      9'd71: begin
        mem_space[71] <= dina;
      end 
      9'd72: begin
        mem_space[72] <= dina;
      end 
      9'd73: begin
        mem_space[73] <= dina;
      end 
      9'd74: begin
        mem_space[74] <= dina;
      end 
      9'd75: begin
        mem_space[75] <= dina;
      end 
      9'd76: begin
        mem_space[76] <= dina;
      end 
      9'd77: begin
        mem_space[77] <= dina;
      end 
      9'd78: begin
        mem_space[78] <= dina;
      end 
      9'd79: begin
        mem_space[79] <= dina;
      end 
      9'd80: begin
        mem_space[80] <= dina;
      end 
      9'd81: begin
        mem_space[81] <= dina;
      end 
      9'd82: begin
        mem_space[82] <= dina;
      end 
      9'd83: begin
        mem_space[83] <= dina;
      end 
      9'd84: begin
        mem_space[84] <= dina;
      end 
      9'd85: begin
        mem_space[85] <= dina;
      end 
      9'd86: begin
        mem_space[86] <= dina;
      end 
      9'd87: begin
        mem_space[87] <= dina;
      end 
      9'd88: begin
        mem_space[88] <= dina;
      end 
      9'd89: begin
        mem_space[89] <= dina;
      end 
      9'd90: begin
        mem_space[90] <= dina;
      end 
      9'd91: begin
        mem_space[91] <= dina;
      end 
      9'd92: begin
        mem_space[92] <= dina;
      end 
      9'd93: begin
        mem_space[93] <= dina;
      end 
      9'd94: begin
        mem_space[94] <= dina;
      end 
      9'd95: begin
        mem_space[95] <= dina;
      end 
      9'd96: begin
        mem_space[96] <= dina;
      end 
      9'd97: begin
        mem_space[97] <= dina;
      end 
      9'd98: begin
        mem_space[98] <= dina;
      end 
      9'd99: begin
        mem_space[99] <= dina;
      end 
      9'd100: begin
        mem_space[100] <= dina;
      end 
      9'd101: begin
        mem_space[101] <= dina;
      end 
      9'd102: begin
        mem_space[102] <= dina;
      end 
      9'd103: begin
        mem_space[103] <= dina;
      end 
      9'd104: begin
        mem_space[104] <= dina;
      end 
      9'd105: begin
        mem_space[105] <= dina;
      end 
      9'd106: begin
        mem_space[106] <= dina;
      end 
      9'd107: begin
        mem_space[107] <= dina;
      end 
      9'd108: begin
        mem_space[108] <= dina;
      end 
      9'd109: begin
        mem_space[109] <= dina;
      end 
      9'd110: begin
        mem_space[110] <= dina;
      end 
      9'd111: begin
        mem_space[111] <= dina;
      end 
      9'd112: begin
        mem_space[112] <= dina;
      end 
      9'd113: begin
        mem_space[113] <= dina;
      end 
      9'd114: begin
        mem_space[114] <= dina;
      end 
      9'd115: begin
        mem_space[115] <= dina;
      end 
      9'd116: begin
        mem_space[116] <= dina;
      end 
      9'd117: begin
        mem_space[117] <= dina;
      end 
      9'd118: begin
        mem_space[118] <= dina;
      end 
      9'd119: begin
        mem_space[119] <= dina;
      end 
      9'd120: begin
        mem_space[120] <= dina;
      end 
      9'd121: begin
        mem_space[121] <= dina;
      end 
      9'd122: begin
        mem_space[122] <= dina;
      end 
      9'd123: begin
        mem_space[123] <= dina;
      end 
      9'd124: begin
        mem_space[124] <= dina;
      end 
      9'd125: begin
        mem_space[125] <= dina;
      end 
      9'd126: begin
        mem_space[126] <= dina;
      end 
      9'd127: begin
        mem_space[127] <= dina;
      end 
      9'd128: begin
        mem_space[128] <= dina;
      end 
      9'd129: begin
        mem_space[129] <= dina;
      end 
      9'd130: begin
        mem_space[130] <= dina;
      end 
      9'd131: begin
        mem_space[131] <= dina;
      end 
      9'd132: begin
        mem_space[132] <= dina;
      end 
      9'd133: begin
        mem_space[133] <= dina;
      end 
      9'd134: begin
        mem_space[134] <= dina;
      end 
      9'd135: begin
        mem_space[135] <= dina;
      end 
      9'd136: begin
        mem_space[136] <= dina;
      end 
      9'd137: begin
        mem_space[137] <= dina;
      end 
      9'd138: begin
        mem_space[138] <= dina;
      end 
      9'd139: begin
        mem_space[139] <= dina;
      end 
      9'd140: begin
        mem_space[140] <= dina;
      end 
      9'd141: begin
        mem_space[141] <= dina;
      end 
      9'd142: begin
        mem_space[142] <= dina;
      end 
      9'd143: begin
        mem_space[143] <= dina;
      end 
      9'd144: begin
        mem_space[144] <= dina;
      end 
      9'd145: begin
        mem_space[145] <= dina;
      end 
      9'd146: begin
        mem_space[146] <= dina;
      end 
      9'd147: begin
        mem_space[147] <= dina;
      end 
      9'd148: begin
        mem_space[148] <= dina;
      end 
      9'd149: begin
        mem_space[149] <= dina;
      end 
      9'd150: begin
        mem_space[150] <= dina;
      end 
      9'd151: begin
        mem_space[151] <= dina;
      end 
      9'd152: begin
        mem_space[152] <= dina;
      end 
      9'd153: begin
        mem_space[153] <= dina;
      end 
      9'd154: begin
        mem_space[154] <= dina;
      end 
      9'd155: begin
        mem_space[155] <= dina;
      end 
      9'd156: begin
        mem_space[156] <= dina;
      end 
      9'd157: begin
        mem_space[157] <= dina;
      end 
      9'd158: begin
        mem_space[158] <= dina;
      end 
      9'd159: begin
        mem_space[159] <= dina;
      end 
      9'd160: begin
        mem_space[160] <= dina;
      end 
      9'd161: begin
        mem_space[161] <= dina;
      end 
      9'd162: begin
        mem_space[162] <= dina;
      end 
      9'd163: begin
        mem_space[163] <= dina;
      end 
      9'd164: begin
        mem_space[164] <= dina;
      end 
      9'd165: begin
        mem_space[165] <= dina;
      end 
      9'd166: begin
        mem_space[166] <= dina;
      end 
      9'd167: begin
        mem_space[167] <= dina;
      end 
      9'd168: begin
        mem_space[168] <= dina;
      end 
      9'd169: begin
        mem_space[169] <= dina;
      end 
      9'd170: begin
        mem_space[170] <= dina;
      end 
      9'd171: begin
        mem_space[171] <= dina;
      end 
      9'd172: begin
        mem_space[172] <= dina;
      end 
      9'd173: begin
        mem_space[173] <= dina;
      end 
      9'd174: begin
        mem_space[174] <= dina;
      end 
      9'd175: begin
        mem_space[175] <= dina;
      end 
      9'd176: begin
        mem_space[176] <= dina;
      end 
      9'd177: begin
        mem_space[177] <= dina;
      end 
      9'd178: begin
        mem_space[178] <= dina;
      end 
      9'd179: begin
        mem_space[179] <= dina;
      end 
      9'd180: begin
        mem_space[180] <= dina;
      end 
      9'd181: begin
        mem_space[181] <= dina;
      end 
      9'd182: begin
        mem_space[182] <= dina;
      end 
      9'd183: begin
        mem_space[183] <= dina;
      end 
      9'd184: begin
        mem_space[184] <= dina;
      end 
      9'd185: begin
        mem_space[185] <= dina;
      end 
      9'd186: begin
        mem_space[186] <= dina;
      end 
      9'd187: begin
        mem_space[187] <= dina;
      end 
      9'd188: begin
        mem_space[188] <= dina;
      end 
      9'd189: begin
        mem_space[189] <= dina;
      end 
      9'd190: begin
        mem_space[190] <= dina;
      end 
      9'd191: begin
        mem_space[191] <= dina;
      end 
      9'd192: begin
        mem_space[192] <= dina;
      end 
      9'd193: begin
        mem_space[193] <= dina;
      end 
      9'd194: begin
        mem_space[194] <= dina;
      end 
      9'd195: begin
        mem_space[195] <= dina;
      end 
      9'd196: begin
        mem_space[196] <= dina;
      end 
      9'd197: begin
        mem_space[197] <= dina;
      end 
      9'd198: begin
        mem_space[198] <= dina;
      end 
      9'd199: begin
        mem_space[199] <= dina;
      end 
      9'd200: begin
        mem_space[200] <= dina;
      end 
      9'd201: begin
        mem_space[201] <= dina;
      end 
      9'd202: begin
        mem_space[202] <= dina;
      end 
      9'd203: begin
        mem_space[203] <= dina;
      end 
      9'd204: begin
        mem_space[204] <= dina;
      end 
      9'd205: begin
        mem_space[205] <= dina;
      end 
      9'd206: begin
        mem_space[206] <= dina;
      end 
      9'd207: begin
        mem_space[207] <= dina;
      end 
      9'd208: begin
        mem_space[208] <= dina;
      end 
      9'd209: begin
        mem_space[209] <= dina;
      end 
      9'd210: begin
        mem_space[210] <= dina;
      end 
      9'd211: begin
        mem_space[211] <= dina;
      end 
      9'd212: begin
        mem_space[212] <= dina;
      end 
      9'd213: begin
        mem_space[213] <= dina;
      end 
      9'd214: begin
        mem_space[214] <= dina;
      end 
      9'd215: begin
        mem_space[215] <= dina;
      end 
      9'd216: begin
        mem_space[216] <= dina;
      end 
      9'd217: begin
        mem_space[217] <= dina;
      end 
      9'd218: begin
        mem_space[218] <= dina;
      end 
      9'd219: begin
        mem_space[219] <= dina;
      end 
      9'd220: begin
        mem_space[220] <= dina;
      end 
      9'd221: begin
        mem_space[221] <= dina;
      end 
      9'd222: begin
        mem_space[222] <= dina;
      end 
      9'd223: begin
        mem_space[223] <= dina;
      end 
      9'd224: begin
        mem_space[224] <= dina;
      end 
      9'd225: begin
        mem_space[225] <= dina;
      end 
      9'd226: begin
        mem_space[226] <= dina;
      end 
      9'd227: begin
        mem_space[227] <= dina;
      end 
      9'd228: begin
        mem_space[228] <= dina;
      end 
      9'd229: begin
        mem_space[229] <= dina;
      end 
      9'd230: begin
        mem_space[230] <= dina;
      end 
      9'd231: begin
        mem_space[231] <= dina;
      end 
      9'd232: begin
        mem_space[232] <= dina;
      end 
      9'd233: begin
        mem_space[233] <= dina;
      end 
      9'd234: begin
        mem_space[234] <= dina;
      end 
      9'd235: begin
        mem_space[235] <= dina;
      end 
      9'd236: begin
        mem_space[236] <= dina;
      end 
      9'd237: begin
        mem_space[237] <= dina;
      end 
      9'd238: begin
        mem_space[238] <= dina;
      end 
      9'd239: begin
        mem_space[239] <= dina;
      end 
      9'd240: begin
        mem_space[240] <= dina;
      end 
      9'd241: begin
        mem_space[241] <= dina;
      end 
      9'd242: begin
        mem_space[242] <= dina;
      end 
      9'd243: begin
        mem_space[243] <= dina;
      end 
      9'd244: begin
        mem_space[244] <= dina;
      end 
      9'd245: begin
        mem_space[245] <= dina;
      end 
      9'd246: begin
        mem_space[246] <= dina;
      end 
      9'd247: begin
        mem_space[247] <= dina;
      end 
      9'd248: begin
        mem_space[248] <= dina;
      end 
      9'd249: begin
        mem_space[249] <= dina;
      end 
      9'd250: begin
        mem_space[250] <= dina;
      end 
      9'd251: begin
        mem_space[251] <= dina;
      end 
      9'd252: begin
        mem_space[252] <= dina;
      end 
      9'd253: begin
        mem_space[253] <= dina;
      end 
      9'd254: begin
        mem_space[254] <= dina;
      end 
      9'd255: begin
        mem_space[255] <= dina;
      end 
      9'd256: begin
        mem_space[256] <= dina;
      end 
      9'd257: begin
        mem_space[257] <= dina;
      end 
      9'd258: begin
        mem_space[258] <= dina;
      end 
      9'd259: begin
        mem_space[259] <= dina;
      end 
      9'd260: begin
        mem_space[260] <= dina;
      end 
      9'd261: begin
        mem_space[261] <= dina;
      end 
      9'd262: begin
        mem_space[262] <= dina;
      end 
      9'd263: begin
        mem_space[263] <= dina;
      end 
      9'd264: begin
        mem_space[264] <= dina;
      end 
      9'd265: begin
        mem_space[265] <= dina;
      end 
      9'd266: begin
        mem_space[266] <= dina;
      end 
      9'd267: begin
        mem_space[267] <= dina;
      end 
      9'd268: begin
        mem_space[268] <= dina;
      end 
      9'd269: begin
        mem_space[269] <= dina;
      end 
      9'd270: begin
        mem_space[270] <= dina;
      end 
      9'd271: begin
        mem_space[271] <= dina;
      end 
      9'd272: begin
        mem_space[272] <= dina;
      end 
      9'd273: begin
        mem_space[273] <= dina;
      end 
      9'd274: begin
        mem_space[274] <= dina;
      end 
      9'd275: begin
        mem_space[275] <= dina;
      end 
      9'd276: begin
        mem_space[276] <= dina;
      end 
      9'd277: begin
        mem_space[277] <= dina;
      end 
      9'd278: begin
        mem_space[278] <= dina;
      end 
      9'd279: begin
        mem_space[279] <= dina;
      end 
      9'd280: begin
        mem_space[280] <= dina;
      end 
      9'd281: begin
        mem_space[281] <= dina;
      end 
      9'd282: begin
        mem_space[282] <= dina;
      end 
      9'd283: begin
        mem_space[283] <= dina;
      end 
      9'd284: begin
        mem_space[284] <= dina;
      end 
      9'd285: begin
        mem_space[285] <= dina;
      end 
      9'd286: begin
        mem_space[286] <= dina;
      end 
      9'd287: begin
        mem_space[287] <= dina;
      end 
      9'd288: begin
        mem_space[288] <= dina;
      end 
      9'd289: begin
        mem_space[289] <= dina;
      end 
      9'd290: begin
        mem_space[290] <= dina;
      end 
      9'd291: begin
        mem_space[291] <= dina;
      end 
      9'd292: begin
        mem_space[292] <= dina;
      end 
      9'd293: begin
        mem_space[293] <= dina;
      end 
      9'd294: begin
        mem_space[294] <= dina;
      end 
      9'd295: begin
        mem_space[295] <= dina;
      end 
      9'd296: begin
        mem_space[296] <= dina;
      end 
      9'd297: begin
        mem_space[297] <= dina;
      end 
      9'd298: begin
        mem_space[298] <= dina;
      end 
      9'd299: begin
        mem_space[299] <= dina;
      end 
      9'd300: begin
        mem_space[300] <= dina;
      end 
      9'd301: begin
        mem_space[301] <= dina;
      end 
      9'd302: begin
        mem_space[302] <= dina;
      end 
      9'd303: begin
        mem_space[303] <= dina;
      end 
      9'd304: begin
        mem_space[304] <= dina;
      end 
      9'd305: begin
        mem_space[305] <= dina;
      end 
      9'd306: begin
        mem_space[306] <= dina;
      end 
      9'd307: begin
        mem_space[307] <= dina;
      end 
      9'd308: begin
        mem_space[308] <= dina;
      end 
      9'd309: begin
        mem_space[309] <= dina;
      end 
      9'd310: begin
        mem_space[310] <= dina;
      end 
      9'd311: begin
        mem_space[311] <= dina;
      end 
      9'd312: begin
        mem_space[312] <= dina;
      end 
      9'd313: begin
        mem_space[313] <= dina;
      end 
      9'd314: begin
        mem_space[314] <= dina;
      end 
      9'd315: begin
        mem_space[315] <= dina;
      end 
      9'd316: begin
        mem_space[316] <= dina;
      end 
      9'd317: begin
        mem_space[317] <= dina;
      end 
      9'd318: begin
        mem_space[318] <= dina;
      end 
      9'd319: begin
        mem_space[319] <= dina;
      end 
      9'd320: begin
        mem_space[320] <= dina;
      end 
      9'd321: begin
        mem_space[321] <= dina;
      end 
      9'd322: begin
        mem_space[322] <= dina;
      end 
      9'd323: begin
        mem_space[323] <= dina;
      end 
      9'd324: begin
        mem_space[324] <= dina;
      end 
      9'd325: begin
        mem_space[325] <= dina;
      end 
      9'd326: begin
        mem_space[326] <= dina;
      end 
      9'd327: begin
        mem_space[327] <= dina;
      end 
      9'd328: begin
        mem_space[328] <= dina;
      end 
      9'd329: begin
        mem_space[329] <= dina;
      end 
      9'd330: begin
        mem_space[330] <= dina;
      end 
      9'd331: begin
        mem_space[331] <= dina;
      end 
      9'd332: begin
        mem_space[332] <= dina;
      end 
      9'd333: begin
        mem_space[333] <= dina;
      end 
      9'd334: begin
        mem_space[334] <= dina;
      end 
      9'd335: begin
        mem_space[335] <= dina;
      end 
      9'd336: begin
        mem_space[336] <= dina;
      end 
      9'd337: begin
        mem_space[337] <= dina;
      end 
      9'd338: begin
        mem_space[338] <= dina;
      end 
      9'd339: begin
        mem_space[339] <= dina;
      end 
      9'd340: begin
        mem_space[340] <= dina;
      end 
      9'd341: begin
        mem_space[341] <= dina;
      end 
      9'd342: begin
        mem_space[342] <= dina;
      end 
      9'd343: begin
        mem_space[343] <= dina;
      end 
      9'd344: begin
        mem_space[344] <= dina;
      end 
      9'd345: begin
        mem_space[345] <= dina;
      end 
      9'd346: begin
        mem_space[346] <= dina;
      end 
      9'd347: begin
        mem_space[347] <= dina;
      end 
      9'd348: begin
        mem_space[348] <= dina;
      end 
      9'd349: begin
        mem_space[349] <= dina;
      end 
      9'd350: begin
        mem_space[350] <= dina;
      end 
      9'd351: begin
        mem_space[351] <= dina;
      end 
      9'd352: begin
        mem_space[352] <= dina;
      end 
      9'd353: begin
        mem_space[353] <= dina;
      end 
      9'd354: begin
        mem_space[354] <= dina;
      end 
      9'd355: begin
        mem_space[355] <= dina;
      end 
      9'd356: begin
        mem_space[356] <= dina;
      end 
      9'd357: begin
        mem_space[357] <= dina;
      end 
      9'd358: begin
        mem_space[358] <= dina;
      end 
      9'd359: begin
        mem_space[359] <= dina;
      end 
      9'd360: begin
        mem_space[360] <= dina;
      end 
      9'd361: begin
        mem_space[361] <= dina;
      end 
      9'd362: begin
        mem_space[362] <= dina;
      end 
      9'd363: begin
        mem_space[363] <= dina;
      end 
      9'd364: begin
        mem_space[364] <= dina;
      end 
      9'd365: begin
        mem_space[365] <= dina;
      end 
      9'd366: begin
        mem_space[366] <= dina;
      end 
      9'd367: begin
        mem_space[367] <= dina;
      end 
      9'd368: begin
        mem_space[368] <= dina;
      end 
      9'd369: begin
        mem_space[369] <= dina;
      end 
      9'd370: begin
        mem_space[370] <= dina;
      end 
      9'd371: begin
        mem_space[371] <= dina;
      end 
      9'd372: begin
        mem_space[372] <= dina;
      end 
      9'd373: begin
        mem_space[373] <= dina;
      end 
      9'd374: begin
        mem_space[374] <= dina;
      end 
      9'd375: begin
        mem_space[375] <= dina;
      end 
      9'd376: begin
        mem_space[376] <= dina;
      end 
      9'd377: begin
        mem_space[377] <= dina;
      end 
      9'd378: begin
        mem_space[378] <= dina;
      end 
      9'd379: begin
        mem_space[379] <= dina;
      end 
      9'd380: begin
        mem_space[380] <= dina;
      end 
      9'd381: begin
        mem_space[381] <= dina;
      end 
      9'd382: begin
        mem_space[382] <= dina;
      end 
      9'd383: begin
        mem_space[383] <= dina;
      end 
      9'd384: begin
        mem_space[384] <= dina;
      end 
      9'd385: begin
        mem_space[385] <= dina;
      end 
      9'd386: begin
        mem_space[386] <= dina;
      end 
      9'd387: begin
        mem_space[387] <= dina;
      end 
      9'd388: begin
        mem_space[388] <= dina;
      end 
      9'd389: begin
        mem_space[389] <= dina;
      end 
      9'd390: begin
        mem_space[390] <= dina;
      end 
      9'd391: begin
        mem_space[391] <= dina;
      end 
      9'd392: begin
        mem_space[392] <= dina;
      end 
      9'd393: begin
        mem_space[393] <= dina;
      end 
      9'd394: begin
        mem_space[394] <= dina;
      end 
      9'd395: begin
        mem_space[395] <= dina;
      end 
      9'd396: begin
        mem_space[396] <= dina;
      end 
      9'd397: begin
        mem_space[397] <= dina;
      end 
      9'd398: begin
        mem_space[398] <= dina;
      end 
      9'd399: begin
        mem_space[399] <= dina;
      end 
      9'd400: begin
        mem_space[400] <= dina;
      end 
      9'd401: begin
        mem_space[401] <= dina;
      end 
      9'd402: begin
        mem_space[402] <= dina;
      end 
      9'd403: begin
        mem_space[403] <= dina;
      end 
      9'd404: begin
        mem_space[404] <= dina;
      end 
      9'd405: begin
        mem_space[405] <= dina;
      end 
      9'd406: begin
        mem_space[406] <= dina;
      end 
      9'd407: begin
        mem_space[407] <= dina;
      end 
      9'd408: begin
        mem_space[408] <= dina;
      end 
      9'd409: begin
        mem_space[409] <= dina;
      end 
      9'd410: begin
        mem_space[410] <= dina;
      end 
      9'd411: begin
        mem_space[411] <= dina;
      end 
      9'd412: begin
        mem_space[412] <= dina;
      end 
      9'd413: begin
        mem_space[413] <= dina;
      end 
      9'd414: begin
        mem_space[414] <= dina;
      end 
      9'd415: begin
        mem_space[415] <= dina;
      end 
      9'd416: begin
        mem_space[416] <= dina;
      end 
      9'd417: begin
        mem_space[417] <= dina;
      end 
      9'd418: begin
        mem_space[418] <= dina;
      end 
      9'd419: begin
        mem_space[419] <= dina;
      end 
      9'd420: begin
        mem_space[420] <= dina;
      end 
      9'd421: begin
        mem_space[421] <= dina;
      end 
      9'd422: begin
        mem_space[422] <= dina;
      end 
      9'd423: begin
        mem_space[423] <= dina;
      end 
      9'd424: begin
        mem_space[424] <= dina;
      end 
      9'd425: begin
        mem_space[425] <= dina;
      end 
      9'd426: begin
        mem_space[426] <= dina;
      end 
      9'd427: begin
        mem_space[427] <= dina;
      end 
      9'd428: begin
        mem_space[428] <= dina;
      end 
      9'd429: begin
        mem_space[429] <= dina;
      end 
      9'd430: begin
        mem_space[430] <= dina;
      end 
      9'd431: begin
        mem_space[431] <= dina;
      end 
      9'd432: begin
        mem_space[432] <= dina;
      end 
      9'd433: begin
        mem_space[433] <= dina;
      end 
      9'd434: begin
        mem_space[434] <= dina;
      end 
      9'd435: begin
        mem_space[435] <= dina;
      end 
      9'd436: begin
        mem_space[436] <= dina;
      end 
      9'd437: begin
        mem_space[437] <= dina;
      end 
      9'd438: begin
        mem_space[438] <= dina;
      end 
      9'd439: begin
        mem_space[439] <= dina;
      end 
      9'd440: begin
        mem_space[440] <= dina;
      end 
      9'd441: begin
        mem_space[441] <= dina;
      end 
      9'd442: begin
        mem_space[442] <= dina;
      end 
      9'd443: begin
        mem_space[443] <= dina;
      end 
      9'd444: begin
        mem_space[444] <= dina;
      end 
      9'd445: begin
        mem_space[445] <= dina;
      end 
      9'd446: begin
        mem_space[446] <= dina;
      end 
      9'd447: begin
        mem_space[447] <= dina;
      end 
      9'd448: begin
        mem_space[448] <= dina;
      end 
      9'd449: begin
        mem_space[449] <= dina;
      end 
      9'd450: begin
        mem_space[450] <= dina;
      end 
      9'd451: begin
        mem_space[451] <= dina;
      end 
      9'd452: begin
        mem_space[452] <= dina;
      end 
      9'd453: begin
        mem_space[453] <= dina;
      end 
      9'd454: begin
        mem_space[454] <= dina;
      end 
      9'd455: begin
        mem_space[455] <= dina;
      end 
      9'd456: begin
        mem_space[456] <= dina;
      end 
      9'd457: begin
        mem_space[457] <= dina;
      end 
      9'd458: begin
        mem_space[458] <= dina;
      end 
      9'd459: begin
        mem_space[459] <= dina;
      end 
      9'd460: begin
        mem_space[460] <= dina;
      end 
      9'd461: begin
        mem_space[461] <= dina;
      end 
      9'd462: begin
        mem_space[462] <= dina;
      end 
      9'd463: begin
        mem_space[463] <= dina;
      end 
      9'd464: begin
        mem_space[464] <= dina;
      end 
      9'd465: begin
        mem_space[465] <= dina;
      end 
      9'd466: begin
        mem_space[466] <= dina;
      end 
      9'd467: begin
        mem_space[467] <= dina;
      end 
      9'd468: begin
        mem_space[468] <= dina;
      end 
      9'd469: begin
        mem_space[469] <= dina;
      end 
      9'd470: begin
        mem_space[470] <= dina;
      end 
      9'd471: begin
        mem_space[471] <= dina;
      end 
      9'd472: begin
        mem_space[472] <= dina;
      end 
      9'd473: begin
        mem_space[473] <= dina;
      end 
      9'd474: begin
        mem_space[474] <= dina;
      end 
      9'd475: begin
        mem_space[475] <= dina;
      end 
      9'd476: begin
        mem_space[476] <= dina;
      end 
      9'd477: begin
        mem_space[477] <= dina;
      end 
      9'd478: begin
        mem_space[478] <= dina;
      end 
      9'd479: begin
        mem_space[479] <= dina;
      end 
      9'd480: begin
        mem_space[480] <= dina;
      end 
      9'd481: begin
        mem_space[481] <= dina;
      end 
      9'd482: begin
        mem_space[482] <= dina;
      end 
      9'd483: begin
        mem_space[483] <= dina;
      end 
      9'd484: begin
        mem_space[484] <= dina;
      end 
      9'd485: begin
        mem_space[485] <= dina;
      end 
      9'd486: begin
        mem_space[486] <= dina;
      end 
      9'd487: begin
        mem_space[487] <= dina;
      end 
      9'd488: begin
        mem_space[488] <= dina;
      end 
      9'd489: begin
        mem_space[489] <= dina;
      end 
      9'd490: begin
        mem_space[490] <= dina;
      end 
      9'd491: begin
        mem_space[491] <= dina;
      end 
      9'd492: begin
        mem_space[492] <= dina;
      end 
      9'd493: begin
        mem_space[493] <= dina;
      end 
      9'd494: begin
        mem_space[494] <= dina;
      end 
      9'd495: begin
        mem_space[495] <= dina;
      end 
      9'd496: begin
        mem_space[496] <= dina;
      end 
      9'd497: begin
        mem_space[497] <= dina;
      end 
      9'd498: begin
        mem_space[498] <= dina;
      end 
      9'd499: begin
        mem_space[499] <= dina;
      end 
      9'd500: begin
        mem_space[500] <= dina;
      end 
      9'd501: begin
        mem_space[501] <= dina;
      end 
      9'd502: begin
        mem_space[502] <= dina;
      end 
      9'd503: begin
        mem_space[503] <= dina;
      end 
      9'd504: begin
        mem_space[504] <= dina;
      end 
      9'd505: begin
        mem_space[505] <= dina;
      end 
      9'd506: begin
        mem_space[506] <= dina;
      end 
      9'd507: begin
        mem_space[507] <= dina;
      end 
      9'd508: begin
        mem_space[508] <= dina;
      end 
      9'd509: begin
        mem_space[509] <= dina;
      end 
      9'd510: begin
        mem_space[510] <= dina;
      end 
      9'd511: begin
        mem_space[511] <= dina;
      end 
      default: begin
        mem_space[0] <= dina;
      end
    endcase
  end
end


always_ff@(posedge clkb) begin
  case ( addr_store ) 
    9'd0: begin
      doutb_pipe <= mem_space[0]; 
    end
    9'd1: begin
      doutb_pipe <= mem_space[1]; 
    end
    9'd2: begin
      doutb_pipe <= mem_space[2]; 
    end
    9'd3: begin
      doutb_pipe <= mem_space[3]; 
    end
    9'd4: begin
      doutb_pipe <= mem_space[4]; 
    end
    9'd5: begin
      doutb_pipe <= mem_space[5]; 
    end
    9'd6: begin
      doutb_pipe <= mem_space[6]; 
    end
    9'd7: begin
      doutb_pipe <= mem_space[7]; 
    end
    9'd8: begin
      doutb_pipe <= mem_space[8]; 
    end
    9'd9: begin
      doutb_pipe <= mem_space[9]; 
    end
    9'd10: begin
      doutb_pipe <= mem_space[10]; 
    end
    9'd11: begin
      doutb_pipe <= mem_space[11]; 
    end
    9'd12: begin
      doutb_pipe <= mem_space[12]; 
    end
    9'd13: begin
      doutb_pipe <= mem_space[13]; 
    end
    9'd14: begin
      doutb_pipe <= mem_space[14]; 
    end
    9'd15: begin
      doutb_pipe <= mem_space[15]; 
    end
    9'd16: begin
      doutb_pipe <= mem_space[16]; 
    end
    9'd17: begin
      doutb_pipe <= mem_space[17]; 
    end
    9'd18: begin
      doutb_pipe <= mem_space[18]; 
    end
    9'd19: begin
      doutb_pipe <= mem_space[19]; 
    end
    9'd20: begin
      doutb_pipe <= mem_space[20]; 
    end
    9'd21: begin
      doutb_pipe <= mem_space[21]; 
    end
    9'd22: begin
      doutb_pipe <= mem_space[22]; 
    end
    9'd23: begin
      doutb_pipe <= mem_space[23]; 
    end
    9'd24: begin
      doutb_pipe <= mem_space[24]; 
    end
    9'd25: begin
      doutb_pipe <= mem_space[25]; 
    end
    9'd26: begin
      doutb_pipe <= mem_space[26]; 
    end
    9'd27: begin
      doutb_pipe <= mem_space[27]; 
    end
    9'd28: begin
      doutb_pipe <= mem_space[28]; 
    end
    9'd29: begin
      doutb_pipe <= mem_space[29]; 
    end
    9'd30: begin
      doutb_pipe <= mem_space[30]; 
    end
    9'd31: begin
      doutb_pipe <= mem_space[31]; 
    end
    9'd32: begin
      doutb_pipe <= mem_space[32]; 
    end
    9'd33: begin
      doutb_pipe <= mem_space[33]; 
    end
    9'd34: begin
      doutb_pipe <= mem_space[34]; 
    end
    9'd35: begin
      doutb_pipe <= mem_space[35]; 
    end
    9'd36: begin
      doutb_pipe <= mem_space[36]; 
    end
    9'd37: begin
      doutb_pipe <= mem_space[37]; 
    end
    9'd38: begin
      doutb_pipe <= mem_space[38]; 
    end
    9'd39: begin
      doutb_pipe <= mem_space[39]; 
    end
    9'd40: begin
      doutb_pipe <= mem_space[40]; 
    end
    9'd41: begin
      doutb_pipe <= mem_space[41]; 
    end
    9'd42: begin
      doutb_pipe <= mem_space[42]; 
    end
    9'd43: begin
      doutb_pipe <= mem_space[43]; 
    end
    9'd44: begin
      doutb_pipe <= mem_space[44]; 
    end
    9'd45: begin
      doutb_pipe <= mem_space[45]; 
    end
    9'd46: begin
      doutb_pipe <= mem_space[46]; 
    end
    9'd47: begin
      doutb_pipe <= mem_space[47]; 
    end
    9'd48: begin
      doutb_pipe <= mem_space[48]; 
    end
    9'd49: begin
      doutb_pipe <= mem_space[49]; 
    end
    9'd50: begin
      doutb_pipe <= mem_space[50]; 
    end
    9'd51: begin
      doutb_pipe <= mem_space[51]; 
    end
    9'd52: begin
      doutb_pipe <= mem_space[52]; 
    end
    9'd53: begin
      doutb_pipe <= mem_space[53]; 
    end
    9'd54: begin
      doutb_pipe <= mem_space[54]; 
    end
    9'd55: begin
      doutb_pipe <= mem_space[55]; 
    end
    9'd56: begin
      doutb_pipe <= mem_space[56]; 
    end
    9'd57: begin
      doutb_pipe <= mem_space[57]; 
    end
    9'd58: begin
      doutb_pipe <= mem_space[58]; 
    end
    9'd59: begin
      doutb_pipe <= mem_space[59]; 
    end
    9'd60: begin
      doutb_pipe <= mem_space[60]; 
    end
    9'd61: begin
      doutb_pipe <= mem_space[61]; 
    end
    9'd62: begin
      doutb_pipe <= mem_space[62]; 
    end
    9'd63: begin
      doutb_pipe <= mem_space[63]; 
    end
    9'd64: begin
      doutb_pipe <= mem_space[64]; 
    end
    9'd65: begin
      doutb_pipe <= mem_space[65]; 
    end
    9'd66: begin
      doutb_pipe <= mem_space[66]; 
    end
    9'd67: begin
      doutb_pipe <= mem_space[67]; 
    end
    9'd68: begin
      doutb_pipe <= mem_space[68]; 
    end
    9'd69: begin
      doutb_pipe <= mem_space[69]; 
    end
    9'd70: begin
      doutb_pipe <= mem_space[70]; 
    end
    9'd71: begin
      doutb_pipe <= mem_space[71]; 
    end
    9'd72: begin
      doutb_pipe <= mem_space[72]; 
    end
    9'd73: begin
      doutb_pipe <= mem_space[73]; 
    end
    9'd74: begin
      doutb_pipe <= mem_space[74]; 
    end
    9'd75: begin
      doutb_pipe <= mem_space[75]; 
    end
    9'd76: begin
      doutb_pipe <= mem_space[76]; 
    end
    9'd77: begin
      doutb_pipe <= mem_space[77]; 
    end
    9'd78: begin
      doutb_pipe <= mem_space[78]; 
    end
    9'd79: begin
      doutb_pipe <= mem_space[79]; 
    end
    9'd80: begin
      doutb_pipe <= mem_space[80]; 
    end
    9'd81: begin
      doutb_pipe <= mem_space[81]; 
    end
    9'd82: begin
      doutb_pipe <= mem_space[82]; 
    end
    9'd83: begin
      doutb_pipe <= mem_space[83]; 
    end
    9'd84: begin
      doutb_pipe <= mem_space[84]; 
    end
    9'd85: begin
      doutb_pipe <= mem_space[85]; 
    end
    9'd86: begin
      doutb_pipe <= mem_space[86]; 
    end
    9'd87: begin
      doutb_pipe <= mem_space[87]; 
    end
    9'd88: begin
      doutb_pipe <= mem_space[88]; 
    end
    9'd89: begin
      doutb_pipe <= mem_space[89]; 
    end
    9'd90: begin
      doutb_pipe <= mem_space[90]; 
    end
    9'd91: begin
      doutb_pipe <= mem_space[91]; 
    end
    9'd92: begin
      doutb_pipe <= mem_space[92]; 
    end
    9'd93: begin
      doutb_pipe <= mem_space[93]; 
    end
    9'd94: begin
      doutb_pipe <= mem_space[94]; 
    end
    9'd95: begin
      doutb_pipe <= mem_space[95]; 
    end
    9'd96: begin
      doutb_pipe <= mem_space[96]; 
    end
    9'd97: begin
      doutb_pipe <= mem_space[97]; 
    end
    9'd98: begin
      doutb_pipe <= mem_space[98]; 
    end
    9'd99: begin
      doutb_pipe <= mem_space[99]; 
    end
    9'd100: begin
      doutb_pipe <= mem_space[100]; 
    end
    9'd101: begin
      doutb_pipe <= mem_space[101]; 
    end
    9'd102: begin
      doutb_pipe <= mem_space[102]; 
    end
    9'd103: begin
      doutb_pipe <= mem_space[103]; 
    end
    9'd104: begin
      doutb_pipe <= mem_space[104]; 
    end
    9'd105: begin
      doutb_pipe <= mem_space[105]; 
    end
    9'd106: begin
      doutb_pipe <= mem_space[106]; 
    end
    9'd107: begin
      doutb_pipe <= mem_space[107]; 
    end
    9'd108: begin
      doutb_pipe <= mem_space[108]; 
    end
    9'd109: begin
      doutb_pipe <= mem_space[109]; 
    end
    9'd110: begin
      doutb_pipe <= mem_space[110]; 
    end
    9'd111: begin
      doutb_pipe <= mem_space[111]; 
    end
    9'd112: begin
      doutb_pipe <= mem_space[112]; 
    end
    9'd113: begin
      doutb_pipe <= mem_space[113]; 
    end
    9'd114: begin
      doutb_pipe <= mem_space[114]; 
    end
    9'd115: begin
      doutb_pipe <= mem_space[115]; 
    end
    9'd116: begin
      doutb_pipe <= mem_space[116]; 
    end
    9'd117: begin
      doutb_pipe <= mem_space[117]; 
    end
    9'd118: begin
      doutb_pipe <= mem_space[118]; 
    end
    9'd119: begin
      doutb_pipe <= mem_space[119]; 
    end
    9'd120: begin
      doutb_pipe <= mem_space[120]; 
    end
    9'd121: begin
      doutb_pipe <= mem_space[121]; 
    end
    9'd122: begin
      doutb_pipe <= mem_space[122]; 
    end
    9'd123: begin
      doutb_pipe <= mem_space[123]; 
    end
    9'd124: begin
      doutb_pipe <= mem_space[124]; 
    end
    9'd125: begin
      doutb_pipe <= mem_space[125]; 
    end
    9'd126: begin
      doutb_pipe <= mem_space[126]; 
    end
    9'd127: begin
      doutb_pipe <= mem_space[127]; 
    end
    9'd128: begin
      doutb_pipe <= mem_space[128]; 
    end
    9'd129: begin
      doutb_pipe <= mem_space[129]; 
    end
    9'd130: begin
      doutb_pipe <= mem_space[130]; 
    end
    9'd131: begin
      doutb_pipe <= mem_space[131]; 
    end
    9'd132: begin
      doutb_pipe <= mem_space[132]; 
    end
    9'd133: begin
      doutb_pipe <= mem_space[133]; 
    end
    9'd134: begin
      doutb_pipe <= mem_space[134]; 
    end
    9'd135: begin
      doutb_pipe <= mem_space[135]; 
    end
    9'd136: begin
      doutb_pipe <= mem_space[136]; 
    end
    9'd137: begin
      doutb_pipe <= mem_space[137]; 
    end
    9'd138: begin
      doutb_pipe <= mem_space[138]; 
    end
    9'd139: begin
      doutb_pipe <= mem_space[139]; 
    end
    9'd140: begin
      doutb_pipe <= mem_space[140]; 
    end
    9'd141: begin
      doutb_pipe <= mem_space[141]; 
    end
    9'd142: begin
      doutb_pipe <= mem_space[142]; 
    end
    9'd143: begin
      doutb_pipe <= mem_space[143]; 
    end
    9'd144: begin
      doutb_pipe <= mem_space[144]; 
    end
    9'd145: begin
      doutb_pipe <= mem_space[145]; 
    end
    9'd146: begin
      doutb_pipe <= mem_space[146]; 
    end
    9'd147: begin
      doutb_pipe <= mem_space[147]; 
    end
    9'd148: begin
      doutb_pipe <= mem_space[148]; 
    end
    9'd149: begin
      doutb_pipe <= mem_space[149]; 
    end
    9'd150: begin
      doutb_pipe <= mem_space[150]; 
    end
    9'd151: begin
      doutb_pipe <= mem_space[151]; 
    end
    9'd152: begin
      doutb_pipe <= mem_space[152]; 
    end
    9'd153: begin
      doutb_pipe <= mem_space[153]; 
    end
    9'd154: begin
      doutb_pipe <= mem_space[154]; 
    end
    9'd155: begin
      doutb_pipe <= mem_space[155]; 
    end
    9'd156: begin
      doutb_pipe <= mem_space[156]; 
    end
    9'd157: begin
      doutb_pipe <= mem_space[157]; 
    end
    9'd158: begin
      doutb_pipe <= mem_space[158]; 
    end
    9'd159: begin
      doutb_pipe <= mem_space[159]; 
    end
    9'd160: begin
      doutb_pipe <= mem_space[160]; 
    end
    9'd161: begin
      doutb_pipe <= mem_space[161]; 
    end
    9'd162: begin
      doutb_pipe <= mem_space[162]; 
    end
    9'd163: begin
      doutb_pipe <= mem_space[163]; 
    end
    9'd164: begin
      doutb_pipe <= mem_space[164]; 
    end
    9'd165: begin
      doutb_pipe <= mem_space[165]; 
    end
    9'd166: begin
      doutb_pipe <= mem_space[166]; 
    end
    9'd167: begin
      doutb_pipe <= mem_space[167]; 
    end
    9'd168: begin
      doutb_pipe <= mem_space[168]; 
    end
    9'd169: begin
      doutb_pipe <= mem_space[169]; 
    end
    9'd170: begin
      doutb_pipe <= mem_space[170]; 
    end
    9'd171: begin
      doutb_pipe <= mem_space[171]; 
    end
    9'd172: begin
      doutb_pipe <= mem_space[172]; 
    end
    9'd173: begin
      doutb_pipe <= mem_space[173]; 
    end
    9'd174: begin
      doutb_pipe <= mem_space[174]; 
    end
    9'd175: begin
      doutb_pipe <= mem_space[175]; 
    end
    9'd176: begin
      doutb_pipe <= mem_space[176]; 
    end
    9'd177: begin
      doutb_pipe <= mem_space[177]; 
    end
    9'd178: begin
      doutb_pipe <= mem_space[178]; 
    end
    9'd179: begin
      doutb_pipe <= mem_space[179]; 
    end
    9'd180: begin
      doutb_pipe <= mem_space[180]; 
    end
    9'd181: begin
      doutb_pipe <= mem_space[181]; 
    end
    9'd182: begin
      doutb_pipe <= mem_space[182]; 
    end
    9'd183: begin
      doutb_pipe <= mem_space[183]; 
    end
    9'd184: begin
      doutb_pipe <= mem_space[184]; 
    end
    9'd185: begin
      doutb_pipe <= mem_space[185]; 
    end
    9'd186: begin
      doutb_pipe <= mem_space[186]; 
    end
    9'd187: begin
      doutb_pipe <= mem_space[187]; 
    end
    9'd188: begin
      doutb_pipe <= mem_space[188]; 
    end
    9'd189: begin
      doutb_pipe <= mem_space[189]; 
    end
    9'd190: begin
      doutb_pipe <= mem_space[190]; 
    end
    9'd191: begin
      doutb_pipe <= mem_space[191]; 
    end
    9'd192: begin
      doutb_pipe <= mem_space[192]; 
    end
    9'd193: begin
      doutb_pipe <= mem_space[193]; 
    end
    9'd194: begin
      doutb_pipe <= mem_space[194]; 
    end
    9'd195: begin
      doutb_pipe <= mem_space[195]; 
    end
    9'd196: begin
      doutb_pipe <= mem_space[196]; 
    end
    9'd197: begin
      doutb_pipe <= mem_space[197]; 
    end
    9'd198: begin
      doutb_pipe <= mem_space[198]; 
    end
    9'd199: begin
      doutb_pipe <= mem_space[199]; 
    end
    9'd200: begin
      doutb_pipe <= mem_space[200]; 
    end
    9'd201: begin
      doutb_pipe <= mem_space[201]; 
    end
    9'd202: begin
      doutb_pipe <= mem_space[202]; 
    end
    9'd203: begin
      doutb_pipe <= mem_space[203]; 
    end
    9'd204: begin
      doutb_pipe <= mem_space[204]; 
    end
    9'd205: begin
      doutb_pipe <= mem_space[205]; 
    end
    9'd206: begin
      doutb_pipe <= mem_space[206]; 
    end
    9'd207: begin
      doutb_pipe <= mem_space[207]; 
    end
    9'd208: begin
      doutb_pipe <= mem_space[208]; 
    end
    9'd209: begin
      doutb_pipe <= mem_space[209]; 
    end
    9'd210: begin
      doutb_pipe <= mem_space[210]; 
    end
    9'd211: begin
      doutb_pipe <= mem_space[211]; 
    end
    9'd212: begin
      doutb_pipe <= mem_space[212]; 
    end
    9'd213: begin
      doutb_pipe <= mem_space[213]; 
    end
    9'd214: begin
      doutb_pipe <= mem_space[214]; 
    end
    9'd215: begin
      doutb_pipe <= mem_space[215]; 
    end
    9'd216: begin
      doutb_pipe <= mem_space[216]; 
    end
    9'd217: begin
      doutb_pipe <= mem_space[217]; 
    end
    9'd218: begin
      doutb_pipe <= mem_space[218]; 
    end
    9'd219: begin
      doutb_pipe <= mem_space[219]; 
    end
    9'd220: begin
      doutb_pipe <= mem_space[220]; 
    end
    9'd221: begin
      doutb_pipe <= mem_space[221]; 
    end
    9'd222: begin
      doutb_pipe <= mem_space[222]; 
    end
    9'd223: begin
      doutb_pipe <= mem_space[223]; 
    end
    9'd224: begin
      doutb_pipe <= mem_space[224]; 
    end
    9'd225: begin
      doutb_pipe <= mem_space[225]; 
    end
    9'd226: begin
      doutb_pipe <= mem_space[226]; 
    end
    9'd227: begin
      doutb_pipe <= mem_space[227]; 
    end
    9'd228: begin
      doutb_pipe <= mem_space[228]; 
    end
    9'd229: begin
      doutb_pipe <= mem_space[229]; 
    end
    9'd230: begin
      doutb_pipe <= mem_space[230]; 
    end
    9'd231: begin
      doutb_pipe <= mem_space[231]; 
    end
    9'd232: begin
      doutb_pipe <= mem_space[232]; 
    end
    9'd233: begin
      doutb_pipe <= mem_space[233]; 
    end
    9'd234: begin
      doutb_pipe <= mem_space[234]; 
    end
    9'd235: begin
      doutb_pipe <= mem_space[235]; 
    end
    9'd236: begin
      doutb_pipe <= mem_space[236]; 
    end
    9'd237: begin
      doutb_pipe <= mem_space[237]; 
    end
    9'd238: begin
      doutb_pipe <= mem_space[238]; 
    end
    9'd239: begin
      doutb_pipe <= mem_space[239]; 
    end
    9'd240: begin
      doutb_pipe <= mem_space[240]; 
    end
    9'd241: begin
      doutb_pipe <= mem_space[241]; 
    end
    9'd242: begin
      doutb_pipe <= mem_space[242]; 
    end
    9'd243: begin
      doutb_pipe <= mem_space[243]; 
    end
    9'd244: begin
      doutb_pipe <= mem_space[244]; 
    end
    9'd245: begin
      doutb_pipe <= mem_space[245]; 
    end
    9'd246: begin
      doutb_pipe <= mem_space[246]; 
    end
    9'd247: begin
      doutb_pipe <= mem_space[247]; 
    end
    9'd248: begin
      doutb_pipe <= mem_space[248]; 
    end
    9'd249: begin
      doutb_pipe <= mem_space[249]; 
    end
    9'd250: begin
      doutb_pipe <= mem_space[250]; 
    end
    9'd251: begin
      doutb_pipe <= mem_space[251]; 
    end
    9'd252: begin
      doutb_pipe <= mem_space[252]; 
    end
    9'd253: begin
      doutb_pipe <= mem_space[253]; 
    end
    9'd254: begin
      doutb_pipe <= mem_space[254]; 
    end
    9'd255: begin
      doutb_pipe <= mem_space[255]; 
    end
    9'd256: begin
      doutb_pipe <= mem_space[256]; 
    end
    9'd257: begin
      doutb_pipe <= mem_space[257]; 
    end
    9'd258: begin
      doutb_pipe <= mem_space[258]; 
    end
    9'd259: begin
      doutb_pipe <= mem_space[259]; 
    end
    9'd260: begin
      doutb_pipe <= mem_space[260]; 
    end
    9'd261: begin
      doutb_pipe <= mem_space[261]; 
    end
    9'd262: begin
      doutb_pipe <= mem_space[262]; 
    end
    9'd263: begin
      doutb_pipe <= mem_space[263]; 
    end
    9'd264: begin
      doutb_pipe <= mem_space[264]; 
    end
    9'd265: begin
      doutb_pipe <= mem_space[265]; 
    end
    9'd266: begin
      doutb_pipe <= mem_space[266]; 
    end
    9'd267: begin
      doutb_pipe <= mem_space[267]; 
    end
    9'd268: begin
      doutb_pipe <= mem_space[268]; 
    end
    9'd269: begin
      doutb_pipe <= mem_space[269]; 
    end
    9'd270: begin
      doutb_pipe <= mem_space[270]; 
    end
    9'd271: begin
      doutb_pipe <= mem_space[271]; 
    end
    9'd272: begin
      doutb_pipe <= mem_space[272]; 
    end
    9'd273: begin
      doutb_pipe <= mem_space[273]; 
    end
    9'd274: begin
      doutb_pipe <= mem_space[274]; 
    end
    9'd275: begin
      doutb_pipe <= mem_space[275]; 
    end
    9'd276: begin
      doutb_pipe <= mem_space[276]; 
    end
    9'd277: begin
      doutb_pipe <= mem_space[277]; 
    end
    9'd278: begin
      doutb_pipe <= mem_space[278]; 
    end
    9'd279: begin
      doutb_pipe <= mem_space[279]; 
    end
    9'd280: begin
      doutb_pipe <= mem_space[280]; 
    end
    9'd281: begin
      doutb_pipe <= mem_space[281]; 
    end
    9'd282: begin
      doutb_pipe <= mem_space[282]; 
    end
    9'd283: begin
      doutb_pipe <= mem_space[283]; 
    end
    9'd284: begin
      doutb_pipe <= mem_space[284]; 
    end
    9'd285: begin
      doutb_pipe <= mem_space[285]; 
    end
    9'd286: begin
      doutb_pipe <= mem_space[286]; 
    end
    9'd287: begin
      doutb_pipe <= mem_space[287]; 
    end
    9'd288: begin
      doutb_pipe <= mem_space[288]; 
    end
    9'd289: begin
      doutb_pipe <= mem_space[289]; 
    end
    9'd290: begin
      doutb_pipe <= mem_space[290]; 
    end
    9'd291: begin
      doutb_pipe <= mem_space[291]; 
    end
    9'd292: begin
      doutb_pipe <= mem_space[292]; 
    end
    9'd293: begin
      doutb_pipe <= mem_space[293]; 
    end
    9'd294: begin
      doutb_pipe <= mem_space[294]; 
    end
    9'd295: begin
      doutb_pipe <= mem_space[295]; 
    end
    9'd296: begin
      doutb_pipe <= mem_space[296]; 
    end
    9'd297: begin
      doutb_pipe <= mem_space[297]; 
    end
    9'd298: begin
      doutb_pipe <= mem_space[298]; 
    end
    9'd299: begin
      doutb_pipe <= mem_space[299]; 
    end
    9'd300: begin
      doutb_pipe <= mem_space[300]; 
    end
    9'd301: begin
      doutb_pipe <= mem_space[301]; 
    end
    9'd302: begin
      doutb_pipe <= mem_space[302]; 
    end
    9'd303: begin
      doutb_pipe <= mem_space[303]; 
    end
    9'd304: begin
      doutb_pipe <= mem_space[304]; 
    end
    9'd305: begin
      doutb_pipe <= mem_space[305]; 
    end
    9'd306: begin
      doutb_pipe <= mem_space[306]; 
    end
    9'd307: begin
      doutb_pipe <= mem_space[307]; 
    end
    9'd308: begin
      doutb_pipe <= mem_space[308]; 
    end
    9'd309: begin
      doutb_pipe <= mem_space[309]; 
    end
    9'd310: begin
      doutb_pipe <= mem_space[310]; 
    end
    9'd311: begin
      doutb_pipe <= mem_space[311]; 
    end
    9'd312: begin
      doutb_pipe <= mem_space[312]; 
    end
    9'd313: begin
      doutb_pipe <= mem_space[313]; 
    end
    9'd314: begin
      doutb_pipe <= mem_space[314]; 
    end
    9'd315: begin
      doutb_pipe <= mem_space[315]; 
    end
    9'd316: begin
      doutb_pipe <= mem_space[316]; 
    end
    9'd317: begin
      doutb_pipe <= mem_space[317]; 
    end
    9'd318: begin
      doutb_pipe <= mem_space[318]; 
    end
    9'd319: begin
      doutb_pipe <= mem_space[319]; 
    end
    9'd320: begin
      doutb_pipe <= mem_space[320]; 
    end
    9'd321: begin
      doutb_pipe <= mem_space[321]; 
    end
    9'd322: begin
      doutb_pipe <= mem_space[322]; 
    end
    9'd323: begin
      doutb_pipe <= mem_space[323]; 
    end
    9'd324: begin
      doutb_pipe <= mem_space[324]; 
    end
    9'd325: begin
      doutb_pipe <= mem_space[325]; 
    end
    9'd326: begin
      doutb_pipe <= mem_space[326]; 
    end
    9'd327: begin
      doutb_pipe <= mem_space[327]; 
    end
    9'd328: begin
      doutb_pipe <= mem_space[328]; 
    end
    9'd329: begin
      doutb_pipe <= mem_space[329]; 
    end
    9'd330: begin
      doutb_pipe <= mem_space[330]; 
    end
    9'd331: begin
      doutb_pipe <= mem_space[331]; 
    end
    9'd332: begin
      doutb_pipe <= mem_space[332]; 
    end
    9'd333: begin
      doutb_pipe <= mem_space[333]; 
    end
    9'd334: begin
      doutb_pipe <= mem_space[334]; 
    end
    9'd335: begin
      doutb_pipe <= mem_space[335]; 
    end
    9'd336: begin
      doutb_pipe <= mem_space[336]; 
    end
    9'd337: begin
      doutb_pipe <= mem_space[337]; 
    end
    9'd338: begin
      doutb_pipe <= mem_space[338]; 
    end
    9'd339: begin
      doutb_pipe <= mem_space[339]; 
    end
    9'd340: begin
      doutb_pipe <= mem_space[340]; 
    end
    9'd341: begin
      doutb_pipe <= mem_space[341]; 
    end
    9'd342: begin
      doutb_pipe <= mem_space[342]; 
    end
    9'd343: begin
      doutb_pipe <= mem_space[343]; 
    end
    9'd344: begin
      doutb_pipe <= mem_space[344]; 
    end
    9'd345: begin
      doutb_pipe <= mem_space[345]; 
    end
    9'd346: begin
      doutb_pipe <= mem_space[346]; 
    end
    9'd347: begin
      doutb_pipe <= mem_space[347]; 
    end
    9'd348: begin
      doutb_pipe <= mem_space[348]; 
    end
    9'd349: begin
      doutb_pipe <= mem_space[349]; 
    end
    9'd350: begin
      doutb_pipe <= mem_space[350]; 
    end
    9'd351: begin
      doutb_pipe <= mem_space[351]; 
    end
    9'd352: begin
      doutb_pipe <= mem_space[352]; 
    end
    9'd353: begin
      doutb_pipe <= mem_space[353]; 
    end
    9'd354: begin
      doutb_pipe <= mem_space[354]; 
    end
    9'd355: begin
      doutb_pipe <= mem_space[355]; 
    end
    9'd356: begin
      doutb_pipe <= mem_space[356]; 
    end
    9'd357: begin
      doutb_pipe <= mem_space[357]; 
    end
    9'd358: begin
      doutb_pipe <= mem_space[358]; 
    end
    9'd359: begin
      doutb_pipe <= mem_space[359]; 
    end
    9'd360: begin
      doutb_pipe <= mem_space[360]; 
    end
    9'd361: begin
      doutb_pipe <= mem_space[361]; 
    end
    9'd362: begin
      doutb_pipe <= mem_space[362]; 
    end
    9'd363: begin
      doutb_pipe <= mem_space[363]; 
    end
    9'd364: begin
      doutb_pipe <= mem_space[364]; 
    end
    9'd365: begin
      doutb_pipe <= mem_space[365]; 
    end
    9'd366: begin
      doutb_pipe <= mem_space[366]; 
    end
    9'd367: begin
      doutb_pipe <= mem_space[367]; 
    end
    9'd368: begin
      doutb_pipe <= mem_space[368]; 
    end
    9'd369: begin
      doutb_pipe <= mem_space[369]; 
    end
    9'd370: begin
      doutb_pipe <= mem_space[370]; 
    end
    9'd371: begin
      doutb_pipe <= mem_space[371]; 
    end
    9'd372: begin
      doutb_pipe <= mem_space[372]; 
    end
    9'd373: begin
      doutb_pipe <= mem_space[373]; 
    end
    9'd374: begin
      doutb_pipe <= mem_space[374]; 
    end
    9'd375: begin
      doutb_pipe <= mem_space[375]; 
    end
    9'd376: begin
      doutb_pipe <= mem_space[376]; 
    end
    9'd377: begin
      doutb_pipe <= mem_space[377]; 
    end
    9'd378: begin
      doutb_pipe <= mem_space[378]; 
    end
    9'd379: begin
      doutb_pipe <= mem_space[379]; 
    end
    9'd380: begin
      doutb_pipe <= mem_space[380]; 
    end
    9'd381: begin
      doutb_pipe <= mem_space[381]; 
    end
    9'd382: begin
      doutb_pipe <= mem_space[382]; 
    end
    9'd383: begin
      doutb_pipe <= mem_space[383]; 
    end
    9'd384: begin
      doutb_pipe <= mem_space[384]; 
    end
    9'd385: begin
      doutb_pipe <= mem_space[385]; 
    end
    9'd386: begin
      doutb_pipe <= mem_space[386]; 
    end
    9'd387: begin
      doutb_pipe <= mem_space[387]; 
    end
    9'd388: begin
      doutb_pipe <= mem_space[388]; 
    end
    9'd389: begin
      doutb_pipe <= mem_space[389]; 
    end
    9'd390: begin
      doutb_pipe <= mem_space[390]; 
    end
    9'd391: begin
      doutb_pipe <= mem_space[391]; 
    end
    9'd392: begin
      doutb_pipe <= mem_space[392]; 
    end
    9'd393: begin
      doutb_pipe <= mem_space[393]; 
    end
    9'd394: begin
      doutb_pipe <= mem_space[394]; 
    end
    9'd395: begin
      doutb_pipe <= mem_space[395]; 
    end
    9'd396: begin
      doutb_pipe <= mem_space[396]; 
    end
    9'd397: begin
      doutb_pipe <= mem_space[397]; 
    end
    9'd398: begin
      doutb_pipe <= mem_space[398]; 
    end
    9'd399: begin
      doutb_pipe <= mem_space[399]; 
    end
    9'd400: begin
      doutb_pipe <= mem_space[400]; 
    end
    9'd401: begin
      doutb_pipe <= mem_space[401]; 
    end
    9'd402: begin
      doutb_pipe <= mem_space[402]; 
    end
    9'd403: begin
      doutb_pipe <= mem_space[403]; 
    end
    9'd404: begin
      doutb_pipe <= mem_space[404]; 
    end
    9'd405: begin
      doutb_pipe <= mem_space[405]; 
    end
    9'd406: begin
      doutb_pipe <= mem_space[406]; 
    end
    9'd407: begin
      doutb_pipe <= mem_space[407]; 
    end
    9'd408: begin
      doutb_pipe <= mem_space[408]; 
    end
    9'd409: begin
      doutb_pipe <= mem_space[409]; 
    end
    9'd410: begin
      doutb_pipe <= mem_space[410]; 
    end
    9'd411: begin
      doutb_pipe <= mem_space[411]; 
    end
    9'd412: begin
      doutb_pipe <= mem_space[412]; 
    end
    9'd413: begin
      doutb_pipe <= mem_space[413]; 
    end
    9'd414: begin
      doutb_pipe <= mem_space[414]; 
    end
    9'd415: begin
      doutb_pipe <= mem_space[415]; 
    end
    9'd416: begin
      doutb_pipe <= mem_space[416]; 
    end
    9'd417: begin
      doutb_pipe <= mem_space[417]; 
    end
    9'd418: begin
      doutb_pipe <= mem_space[418]; 
    end
    9'd419: begin
      doutb_pipe <= mem_space[419]; 
    end
    9'd420: begin
      doutb_pipe <= mem_space[420]; 
    end
    9'd421: begin
      doutb_pipe <= mem_space[421]; 
    end
    9'd422: begin
      doutb_pipe <= mem_space[422]; 
    end
    9'd423: begin
      doutb_pipe <= mem_space[423]; 
    end
    9'd424: begin
      doutb_pipe <= mem_space[424]; 
    end
    9'd425: begin
      doutb_pipe <= mem_space[425]; 
    end
    9'd426: begin
      doutb_pipe <= mem_space[426]; 
    end
    9'd427: begin
      doutb_pipe <= mem_space[427]; 
    end
    9'd428: begin
      doutb_pipe <= mem_space[428]; 
    end
    9'd429: begin
      doutb_pipe <= mem_space[429]; 
    end
    9'd430: begin
      doutb_pipe <= mem_space[430]; 
    end
    9'd431: begin
      doutb_pipe <= mem_space[431]; 
    end
    9'd432: begin
      doutb_pipe <= mem_space[432]; 
    end
    9'd433: begin
      doutb_pipe <= mem_space[433]; 
    end
    9'd434: begin
      doutb_pipe <= mem_space[434]; 
    end
    9'd435: begin
      doutb_pipe <= mem_space[435]; 
    end
    9'd436: begin
      doutb_pipe <= mem_space[436]; 
    end
    9'd437: begin
      doutb_pipe <= mem_space[437]; 
    end
    9'd438: begin
      doutb_pipe <= mem_space[438]; 
    end
    9'd439: begin
      doutb_pipe <= mem_space[439]; 
    end
    9'd440: begin
      doutb_pipe <= mem_space[440]; 
    end
    9'd441: begin
      doutb_pipe <= mem_space[441]; 
    end
    9'd442: begin
      doutb_pipe <= mem_space[442]; 
    end
    9'd443: begin
      doutb_pipe <= mem_space[443]; 
    end
    9'd444: begin
      doutb_pipe <= mem_space[444]; 
    end
    9'd445: begin
      doutb_pipe <= mem_space[445]; 
    end
    9'd446: begin
      doutb_pipe <= mem_space[446]; 
    end
    9'd447: begin
      doutb_pipe <= mem_space[447]; 
    end
    9'd448: begin
      doutb_pipe <= mem_space[448]; 
    end
    9'd449: begin
      doutb_pipe <= mem_space[449]; 
    end
    9'd450: begin
      doutb_pipe <= mem_space[450]; 
    end
    9'd451: begin
      doutb_pipe <= mem_space[451]; 
    end
    9'd452: begin
      doutb_pipe <= mem_space[452]; 
    end
    9'd453: begin
      doutb_pipe <= mem_space[453]; 
    end
    9'd454: begin
      doutb_pipe <= mem_space[454]; 
    end
    9'd455: begin
      doutb_pipe <= mem_space[455]; 
    end
    9'd456: begin
      doutb_pipe <= mem_space[456]; 
    end
    9'd457: begin
      doutb_pipe <= mem_space[457]; 
    end
    9'd458: begin
      doutb_pipe <= mem_space[458]; 
    end
    9'd459: begin
      doutb_pipe <= mem_space[459]; 
    end
    9'd460: begin
      doutb_pipe <= mem_space[460]; 
    end
    9'd461: begin
      doutb_pipe <= mem_space[461]; 
    end
    9'd462: begin
      doutb_pipe <= mem_space[462]; 
    end
    9'd463: begin
      doutb_pipe <= mem_space[463]; 
    end
    9'd464: begin
      doutb_pipe <= mem_space[464]; 
    end
    9'd465: begin
      doutb_pipe <= mem_space[465]; 
    end
    9'd466: begin
      doutb_pipe <= mem_space[466]; 
    end
    9'd467: begin
      doutb_pipe <= mem_space[467]; 
    end
    9'd468: begin
      doutb_pipe <= mem_space[468]; 
    end
    9'd469: begin
      doutb_pipe <= mem_space[469]; 
    end
    9'd470: begin
      doutb_pipe <= mem_space[470]; 
    end
    9'd471: begin
      doutb_pipe <= mem_space[471]; 
    end
    9'd472: begin
      doutb_pipe <= mem_space[472]; 
    end
    9'd473: begin
      doutb_pipe <= mem_space[473]; 
    end
    9'd474: begin
      doutb_pipe <= mem_space[474]; 
    end
    9'd475: begin
      doutb_pipe <= mem_space[475]; 
    end
    9'd476: begin
      doutb_pipe <= mem_space[476]; 
    end
    9'd477: begin
      doutb_pipe <= mem_space[477]; 
    end
    9'd478: begin
      doutb_pipe <= mem_space[478]; 
    end
    9'd479: begin
      doutb_pipe <= mem_space[479]; 
    end
    9'd480: begin
      doutb_pipe <= mem_space[480]; 
    end
    9'd481: begin
      doutb_pipe <= mem_space[481]; 
    end
    9'd482: begin
      doutb_pipe <= mem_space[482]; 
    end
    9'd483: begin
      doutb_pipe <= mem_space[483]; 
    end
    9'd484: begin
      doutb_pipe <= mem_space[484]; 
    end
    9'd485: begin
      doutb_pipe <= mem_space[485]; 
    end
    9'd486: begin
      doutb_pipe <= mem_space[486]; 
    end
    9'd487: begin
      doutb_pipe <= mem_space[487]; 
    end
    9'd488: begin
      doutb_pipe <= mem_space[488]; 
    end
    9'd489: begin
      doutb_pipe <= mem_space[489]; 
    end
    9'd490: begin
      doutb_pipe <= mem_space[490]; 
    end
    9'd491: begin
      doutb_pipe <= mem_space[491]; 
    end
    9'd492: begin
      doutb_pipe <= mem_space[492]; 
    end
    9'd493: begin
      doutb_pipe <= mem_space[493]; 
    end
    9'd494: begin
      doutb_pipe <= mem_space[494]; 
    end
    9'd495: begin
      doutb_pipe <= mem_space[495]; 
    end
    9'd496: begin
      doutb_pipe <= mem_space[496]; 
    end
    9'd497: begin
      doutb_pipe <= mem_space[497]; 
    end
    9'd498: begin
      doutb_pipe <= mem_space[498]; 
    end
    9'd499: begin
      doutb_pipe <= mem_space[499]; 
    end
    9'd500: begin
      doutb_pipe <= mem_space[500]; 
    end
    9'd501: begin
      doutb_pipe <= mem_space[501]; 
    end
    9'd502: begin
      doutb_pipe <= mem_space[502]; 
    end
    9'd503: begin
      doutb_pipe <= mem_space[503]; 
    end
    9'd504: begin
      doutb_pipe <= mem_space[504]; 
    end
    9'd505: begin
      doutb_pipe <= mem_space[505]; 
    end
    9'd506: begin
      doutb_pipe <= mem_space[506]; 
    end
    9'd507: begin
      doutb_pipe <= mem_space[507]; 
    end
    9'd508: begin
      doutb_pipe <= mem_space[508]; 
    end
    9'd509: begin
      doutb_pipe <= mem_space[509]; 
    end
    9'd510: begin
      doutb_pipe <= mem_space[510]; 
    end
    9'd511: begin
      doutb_pipe <= mem_space[511]; 
    end
    default: begin
      doutb_pipe <= '0;
    end
  endcase
end

always_ff@(posedge clkb) begin
  if ( enb ) begin
    addr_store <= addrb;
  end
end

always_ff@(posedge clkb) begin
  doutb <= doutb_pipe;
end



endmodule
