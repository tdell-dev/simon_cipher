module simon_fifo (
  input wire clk,
  input wire srst,

  input wire [7:0] din,
  input wire wr_en,

  output logic [7:0] dout,
  input wire rd_en,

  output logic empty,
  output logic full,

  output logic wr_rst_busy,
  output logic rd_rst_busy
);

//There are 512 entries, expand it out

logic [8:0] waddr;
logic [8:0] raddr;
logic [511:0][7:0] mem_space;

assign empty = waddr == raddr;
assign full = waddr+1 == raddr;

always_ff@(posedge clk) begin
  if ( srst ) begin
    waddr <= '0;
    raddr <= '0;
  end
end

always_ff@(posedge clk) begin
  if ( wr_en ) begin
    waddr <= waddr + 1;
  end
end

always_ff@(posedge clk) begin
  if ( rd_en ) begin
    raddr <= raddr + 1;
  end
end

always_ff@(posedge clk) begin
  case( raddr )
    9'd0: begin
      dout <= mem_space[0];
    end
    9'd1: begin
      dout <= mem_space[1];
    end
    9'd2: begin
      dout <= mem_space[2];
    end
    9'd3: begin
      dout <= mem_space[3];
    end
    9'd4: begin
      dout <= mem_space[4];
    end
    9'd5: begin
      dout <= mem_space[5];
    end
    9'd6: begin
      dout <= mem_space[6];
    end
    9'd7: begin
      dout <= mem_space[7];
    end
    9'd8: begin
      dout <= mem_space[8];
    end
    9'd9: begin
      dout <= mem_space[9];
    end
    9'd10: begin
      dout <= mem_space[10];
    end
    9'd11: begin
      dout <= mem_space[11];
    end
    9'd12: begin
      dout <= mem_space[12];
    end
    9'd13: begin
      dout <= mem_space[13];
    end
    9'd14: begin
      dout <= mem_space[14];
    end
    9'd15: begin
      dout <= mem_space[15];
    end
    9'd16: begin
      dout <= mem_space[16];
    end
    9'd17: begin
      dout <= mem_space[17];
    end
    9'd18: begin
      dout <= mem_space[18];
    end
    9'd19: begin
      dout <= mem_space[19];
    end
    9'd20: begin
      dout <= mem_space[20];
    end
    9'd21: begin
      dout <= mem_space[21];
    end
    9'd22: begin
      dout <= mem_space[22];
    end
    9'd23: begin
      dout <= mem_space[23];
    end
    9'd24: begin
      dout <= mem_space[24];
    end
    9'd25: begin
      dout <= mem_space[25];
    end
    9'd26: begin
      dout <= mem_space[26];
    end
    9'd27: begin
      dout <= mem_space[27];
    end
    9'd28: begin
      dout <= mem_space[28];
    end
    9'd29: begin
      dout <= mem_space[29];
    end
    9'd30: begin
      dout <= mem_space[30];
    end
    9'd31: begin
      dout <= mem_space[31];
    end
    9'd32: begin
      dout <= mem_space[32];
    end
    9'd33: begin
      dout <= mem_space[33];
    end
    9'd34: begin
      dout <= mem_space[34];
    end
    9'd35: begin
      dout <= mem_space[35];
    end
    9'd36: begin
      dout <= mem_space[36];
    end
    9'd37: begin
      dout <= mem_space[37];
    end
    9'd38: begin
      dout <= mem_space[38];
    end
    9'd39: begin
      dout <= mem_space[39];
    end
    9'd40: begin
      dout <= mem_space[40];
    end
    9'd41: begin
      dout <= mem_space[41];
    end
    9'd42: begin
      dout <= mem_space[42];
    end
    9'd43: begin
      dout <= mem_space[43];
    end
    9'd44: begin
      dout <= mem_space[44];
    end
    9'd45: begin
      dout <= mem_space[45];
    end
    9'd46: begin
      dout <= mem_space[46];
    end
    9'd47: begin
      dout <= mem_space[47];
    end
    9'd48: begin
      dout <= mem_space[48];
    end
    9'd49: begin
      dout <= mem_space[49];
    end
    9'd50: begin
      dout <= mem_space[50];
    end
    9'd51: begin
      dout <= mem_space[51];
    end
    9'd52: begin
      dout <= mem_space[52];
    end
    9'd53: begin
      dout <= mem_space[53];
    end
    9'd54: begin
      dout <= mem_space[54];
    end
    9'd55: begin
      dout <= mem_space[55];
    end
    9'd56: begin
      dout <= mem_space[56];
    end
    9'd57: begin
      dout <= mem_space[57];
    end
    9'd58: begin
      dout <= mem_space[58];
    end
    9'd59: begin
      dout <= mem_space[59];
    end
    9'd60: begin
      dout <= mem_space[60];
    end
    9'd61: begin
      dout <= mem_space[61];
    end
    9'd62: begin
      dout <= mem_space[62];
    end
    9'd63: begin
      dout <= mem_space[63];
    end
    9'd64: begin
      dout <= mem_space[64];
    end
    9'd65: begin
      dout <= mem_space[65];
    end
    9'd66: begin
      dout <= mem_space[66];
    end
    9'd67: begin
      dout <= mem_space[67];
    end
    9'd68: begin
      dout <= mem_space[68];
    end
    9'd69: begin
      dout <= mem_space[69];
    end
    9'd70: begin
      dout <= mem_space[70];
    end
    9'd71: begin
      dout <= mem_space[71];
    end
    9'd72: begin
      dout <= mem_space[72];
    end
    9'd73: begin
      dout <= mem_space[73];
    end
    9'd74: begin
      dout <= mem_space[74];
    end
    9'd75: begin
      dout <= mem_space[75];
    end
    9'd76: begin
      dout <= mem_space[76];
    end
    9'd77: begin
      dout <= mem_space[77];
    end
    9'd78: begin
      dout <= mem_space[78];
    end
    9'd79: begin
      dout <= mem_space[79];
    end
    9'd80: begin
      dout <= mem_space[80];
    end
    9'd81: begin
      dout <= mem_space[81];
    end
    9'd82: begin
      dout <= mem_space[82];
    end
    9'd83: begin
      dout <= mem_space[83];
    end
    9'd84: begin
      dout <= mem_space[84];
    end
    9'd85: begin
      dout <= mem_space[85];
    end
    9'd86: begin
      dout <= mem_space[86];
    end
    9'd87: begin
      dout <= mem_space[87];
    end
    9'd88: begin
      dout <= mem_space[88];
    end
    9'd89: begin
      dout <= mem_space[89];
    end
    9'd90: begin
      dout <= mem_space[90];
    end
    9'd91: begin
      dout <= mem_space[91];
    end
    9'd92: begin
      dout <= mem_space[92];
    end
    9'd93: begin
      dout <= mem_space[93];
    end
    9'd94: begin
      dout <= mem_space[94];
    end
    9'd95: begin
      dout <= mem_space[95];
    end
    9'd96: begin
      dout <= mem_space[96];
    end
    9'd97: begin
      dout <= mem_space[97];
    end
    9'd98: begin
      dout <= mem_space[98];
    end
    9'd99: begin
      dout <= mem_space[99];
    end
    9'd100: begin
      dout <= mem_space[100];
    end
    9'd101: begin
      dout <= mem_space[101];
    end
    9'd102: begin
      dout <= mem_space[102];
    end
    9'd103: begin
      dout <= mem_space[103];
    end
    9'd104: begin
      dout <= mem_space[104];
    end
    9'd105: begin
      dout <= mem_space[105];
    end
    9'd106: begin
      dout <= mem_space[106];
    end
    9'd107: begin
      dout <= mem_space[107];
    end
    9'd108: begin
      dout <= mem_space[108];
    end
    9'd109: begin
      dout <= mem_space[109];
    end
    9'd110: begin
      dout <= mem_space[110];
    end
    9'd111: begin
      dout <= mem_space[111];
    end
    9'd112: begin
      dout <= mem_space[112];
    end
    9'd113: begin
      dout <= mem_space[113];
    end
    9'd114: begin
      dout <= mem_space[114];
    end
    9'd115: begin
      dout <= mem_space[115];
    end
    9'd116: begin
      dout <= mem_space[116];
    end
    9'd117: begin
      dout <= mem_space[117];
    end
    9'd118: begin
      dout <= mem_space[118];
    end
    9'd119: begin
      dout <= mem_space[119];
    end
    9'd120: begin
      dout <= mem_space[120];
    end
    9'd121: begin
      dout <= mem_space[121];
    end
    9'd122: begin
      dout <= mem_space[122];
    end
    9'd123: begin
      dout <= mem_space[123];
    end
    9'd124: begin
      dout <= mem_space[124];
    end
    9'd125: begin
      dout <= mem_space[125];
    end
    9'd126: begin
      dout <= mem_space[126];
    end
    9'd127: begin
      dout <= mem_space[127];
    end
    9'd128: begin
      dout <= mem_space[128];
    end
    9'd129: begin
      dout <= mem_space[129];
    end
    9'd130: begin
      dout <= mem_space[130];
    end
    9'd131: begin
      dout <= mem_space[131];
    end
    9'd132: begin
      dout <= mem_space[132];
    end
    9'd133: begin
      dout <= mem_space[133];
    end
    9'd134: begin
      dout <= mem_space[134];
    end
    9'd135: begin
      dout <= mem_space[135];
    end
    9'd136: begin
      dout <= mem_space[136];
    end
    9'd137: begin
      dout <= mem_space[137];
    end
    9'd138: begin
      dout <= mem_space[138];
    end
    9'd139: begin
      dout <= mem_space[139];
    end
    9'd140: begin
      dout <= mem_space[140];
    end
    9'd141: begin
      dout <= mem_space[141];
    end
    9'd142: begin
      dout <= mem_space[142];
    end
    9'd143: begin
      dout <= mem_space[143];
    end
    9'd144: begin
      dout <= mem_space[144];
    end
    9'd145: begin
      dout <= mem_space[145];
    end
    9'd146: begin
      dout <= mem_space[146];
    end
    9'd147: begin
      dout <= mem_space[147];
    end
    9'd148: begin
      dout <= mem_space[148];
    end
    9'd149: begin
      dout <= mem_space[149];
    end
    9'd150: begin
      dout <= mem_space[150];
    end
    9'd151: begin
      dout <= mem_space[151];
    end
    9'd152: begin
      dout <= mem_space[152];
    end
    9'd153: begin
      dout <= mem_space[153];
    end
    9'd154: begin
      dout <= mem_space[154];
    end
    9'd155: begin
      dout <= mem_space[155];
    end
    9'd156: begin
      dout <= mem_space[156];
    end
    9'd157: begin
      dout <= mem_space[157];
    end
    9'd158: begin
      dout <= mem_space[158];
    end
    9'd159: begin
      dout <= mem_space[159];
    end
    9'd160: begin
      dout <= mem_space[160];
    end
    9'd161: begin
      dout <= mem_space[161];
    end
    9'd162: begin
      dout <= mem_space[162];
    end
    9'd163: begin
      dout <= mem_space[163];
    end
    9'd164: begin
      dout <= mem_space[164];
    end
    9'd165: begin
      dout <= mem_space[165];
    end
    9'd166: begin
      dout <= mem_space[166];
    end
    9'd167: begin
      dout <= mem_space[167];
    end
    9'd168: begin
      dout <= mem_space[168];
    end
    9'd169: begin
      dout <= mem_space[169];
    end
    9'd170: begin
      dout <= mem_space[170];
    end
    9'd171: begin
      dout <= mem_space[171];
    end
    9'd172: begin
      dout <= mem_space[172];
    end
    9'd173: begin
      dout <= mem_space[173];
    end
    9'd174: begin
      dout <= mem_space[174];
    end
    9'd175: begin
      dout <= mem_space[175];
    end
    9'd176: begin
      dout <= mem_space[176];
    end
    9'd177: begin
      dout <= mem_space[177];
    end
    9'd178: begin
      dout <= mem_space[178];
    end
    9'd179: begin
      dout <= mem_space[179];
    end
    9'd180: begin
      dout <= mem_space[180];
    end
    9'd181: begin
      dout <= mem_space[181];
    end
    9'd182: begin
      dout <= mem_space[182];
    end
    9'd183: begin
      dout <= mem_space[183];
    end
    9'd184: begin
      dout <= mem_space[184];
    end
    9'd185: begin
      dout <= mem_space[185];
    end
    9'd186: begin
      dout <= mem_space[186];
    end
    9'd187: begin
      dout <= mem_space[187];
    end
    9'd188: begin
      dout <= mem_space[188];
    end
    9'd189: begin
      dout <= mem_space[189];
    end
    9'd190: begin
      dout <= mem_space[190];
    end
    9'd191: begin
      dout <= mem_space[191];
    end
    9'd192: begin
      dout <= mem_space[192];
    end
    9'd193: begin
      dout <= mem_space[193];
    end
    9'd194: begin
      dout <= mem_space[194];
    end
    9'd195: begin
      dout <= mem_space[195];
    end
    9'd196: begin
      dout <= mem_space[196];
    end
    9'd197: begin
      dout <= mem_space[197];
    end
    9'd198: begin
      dout <= mem_space[198];
    end
    9'd199: begin
      dout <= mem_space[199];
    end
    9'd200: begin
      dout <= mem_space[200];
    end
    9'd201: begin
      dout <= mem_space[201];
    end
    9'd202: begin
      dout <= mem_space[202];
    end
    9'd203: begin
      dout <= mem_space[203];
    end
    9'd204: begin
      dout <= mem_space[204];
    end
    9'd205: begin
      dout <= mem_space[205];
    end
    9'd206: begin
      dout <= mem_space[206];
    end
    9'd207: begin
      dout <= mem_space[207];
    end
    9'd208: begin
      dout <= mem_space[208];
    end
    9'd209: begin
      dout <= mem_space[209];
    end
    9'd210: begin
      dout <= mem_space[210];
    end
    9'd211: begin
      dout <= mem_space[211];
    end
    9'd212: begin
      dout <= mem_space[212];
    end
    9'd213: begin
      dout <= mem_space[213];
    end
    9'd214: begin
      dout <= mem_space[214];
    end
    9'd215: begin
      dout <= mem_space[215];
    end
    9'd216: begin
      dout <= mem_space[216];
    end
    9'd217: begin
      dout <= mem_space[217];
    end
    9'd218: begin
      dout <= mem_space[218];
    end
    9'd219: begin
      dout <= mem_space[219];
    end
    9'd220: begin
      dout <= mem_space[220];
    end
    9'd221: begin
      dout <= mem_space[221];
    end
    9'd222: begin
      dout <= mem_space[222];
    end
    9'd223: begin
      dout <= mem_space[223];
    end
    9'd224: begin
      dout <= mem_space[224];
    end
    9'd225: begin
      dout <= mem_space[225];
    end
    9'd226: begin
      dout <= mem_space[226];
    end
    9'd227: begin
      dout <= mem_space[227];
    end
    9'd228: begin
      dout <= mem_space[228];
    end
    9'd229: begin
      dout <= mem_space[229];
    end
    9'd230: begin
      dout <= mem_space[230];
    end
    9'd231: begin
      dout <= mem_space[231];
    end
    9'd232: begin
      dout <= mem_space[232];
    end
    9'd233: begin
      dout <= mem_space[233];
    end
    9'd234: begin
      dout <= mem_space[234];
    end
    9'd235: begin
      dout <= mem_space[235];
    end
    9'd236: begin
      dout <= mem_space[236];
    end
    9'd237: begin
      dout <= mem_space[237];
    end
    9'd238: begin
      dout <= mem_space[238];
    end
    9'd239: begin
      dout <= mem_space[239];
    end
    9'd240: begin
      dout <= mem_space[240];
    end
    9'd241: begin
      dout <= mem_space[241];
    end
    9'd242: begin
      dout <= mem_space[242];
    end
    9'd243: begin
      dout <= mem_space[243];
    end
    9'd244: begin
      dout <= mem_space[244];
    end
    9'd245: begin
      dout <= mem_space[245];
    end
    9'd246: begin
      dout <= mem_space[246];
    end
    9'd247: begin
      dout <= mem_space[247];
    end
    9'd248: begin
      dout <= mem_space[248];
    end
    9'd249: begin
      dout <= mem_space[249];
    end
    9'd250: begin
      dout <= mem_space[250];
    end
    9'd251: begin
      dout <= mem_space[251];
    end
    9'd252: begin
      dout <= mem_space[252];
    end
    9'd253: begin
      dout <= mem_space[253];
    end
    9'd254: begin
      dout <= mem_space[254];
    end
    9'd255: begin
      dout <= mem_space[255];
    end
    9'd256: begin
      dout <= mem_space[256];
    end
    9'd257: begin
      dout <= mem_space[257];
    end
    9'd258: begin
      dout <= mem_space[258];
    end
    9'd259: begin
      dout <= mem_space[259];
    end
    9'd260: begin
      dout <= mem_space[260];
    end
    9'd261: begin
      dout <= mem_space[261];
    end
    9'd262: begin
      dout <= mem_space[262];
    end
    9'd263: begin
      dout <= mem_space[263];
    end
    9'd264: begin
      dout <= mem_space[264];
    end
    9'd265: begin
      dout <= mem_space[265];
    end
    9'd266: begin
      dout <= mem_space[266];
    end
    9'd267: begin
      dout <= mem_space[267];
    end
    9'd268: begin
      dout <= mem_space[268];
    end
    9'd269: begin
      dout <= mem_space[269];
    end
    9'd270: begin
      dout <= mem_space[270];
    end
    9'd271: begin
      dout <= mem_space[271];
    end
    9'd272: begin
      dout <= mem_space[272];
    end
    9'd273: begin
      dout <= mem_space[273];
    end
    9'd274: begin
      dout <= mem_space[274];
    end
    9'd275: begin
      dout <= mem_space[275];
    end
    9'd276: begin
      dout <= mem_space[276];
    end
    9'd277: begin
      dout <= mem_space[277];
    end
    9'd278: begin
      dout <= mem_space[278];
    end
    9'd279: begin
      dout <= mem_space[279];
    end
    9'd280: begin
      dout <= mem_space[280];
    end
    9'd281: begin
      dout <= mem_space[281];
    end
    9'd282: begin
      dout <= mem_space[282];
    end
    9'd283: begin
      dout <= mem_space[283];
    end
    9'd284: begin
      dout <= mem_space[284];
    end
    9'd285: begin
      dout <= mem_space[285];
    end
    9'd286: begin
      dout <= mem_space[286];
    end
    9'd287: begin
      dout <= mem_space[287];
    end
    9'd288: begin
      dout <= mem_space[288];
    end
    9'd289: begin
      dout <= mem_space[289];
    end
    9'd290: begin
      dout <= mem_space[290];
    end
    9'd291: begin
      dout <= mem_space[291];
    end
    9'd292: begin
      dout <= mem_space[292];
    end
    9'd293: begin
      dout <= mem_space[293];
    end
    9'd294: begin
      dout <= mem_space[294];
    end
    9'd295: begin
      dout <= mem_space[295];
    end
    9'd296: begin
      dout <= mem_space[296];
    end
    9'd297: begin
      dout <= mem_space[297];
    end
    9'd298: begin
      dout <= mem_space[298];
    end
    9'd299: begin
      dout <= mem_space[299];
    end
    9'd300: begin
      dout <= mem_space[300];
    end
    9'd301: begin
      dout <= mem_space[301];
    end
    9'd302: begin
      dout <= mem_space[302];
    end
    9'd303: begin
      dout <= mem_space[303];
    end
    9'd304: begin
      dout <= mem_space[304];
    end
    9'd305: begin
      dout <= mem_space[305];
    end
    9'd306: begin
      dout <= mem_space[306];
    end
    9'd307: begin
      dout <= mem_space[307];
    end
    9'd308: begin
      dout <= mem_space[308];
    end
    9'd309: begin
      dout <= mem_space[309];
    end
    9'd310: begin
      dout <= mem_space[310];
    end
    9'd311: begin
      dout <= mem_space[311];
    end
    9'd312: begin
      dout <= mem_space[312];
    end
    9'd313: begin
      dout <= mem_space[313];
    end
    9'd314: begin
      dout <= mem_space[314];
    end
    9'd315: begin
      dout <= mem_space[315];
    end
    9'd316: begin
      dout <= mem_space[316];
    end
    9'd317: begin
      dout <= mem_space[317];
    end
    9'd318: begin
      dout <= mem_space[318];
    end
    9'd319: begin
      dout <= mem_space[319];
    end
    9'd320: begin
      dout <= mem_space[320];
    end
    9'd321: begin
      dout <= mem_space[321];
    end
    9'd322: begin
      dout <= mem_space[322];
    end
    9'd323: begin
      dout <= mem_space[323];
    end
    9'd324: begin
      dout <= mem_space[324];
    end
    9'd325: begin
      dout <= mem_space[325];
    end
    9'd326: begin
      dout <= mem_space[326];
    end
    9'd327: begin
      dout <= mem_space[327];
    end
    9'd328: begin
      dout <= mem_space[328];
    end
    9'd329: begin
      dout <= mem_space[329];
    end
    9'd330: begin
      dout <= mem_space[330];
    end
    9'd331: begin
      dout <= mem_space[331];
    end
    9'd332: begin
      dout <= mem_space[332];
    end
    9'd333: begin
      dout <= mem_space[333];
    end
    9'd334: begin
      dout <= mem_space[334];
    end
    9'd335: begin
      dout <= mem_space[335];
    end
    9'd336: begin
      dout <= mem_space[336];
    end
    9'd337: begin
      dout <= mem_space[337];
    end
    9'd338: begin
      dout <= mem_space[338];
    end
    9'd339: begin
      dout <= mem_space[339];
    end
    9'd340: begin
      dout <= mem_space[340];
    end
    9'd341: begin
      dout <= mem_space[341];
    end
    9'd342: begin
      dout <= mem_space[342];
    end
    9'd343: begin
      dout <= mem_space[343];
    end
    9'd344: begin
      dout <= mem_space[344];
    end
    9'd345: begin
      dout <= mem_space[345];
    end
    9'd346: begin
      dout <= mem_space[346];
    end
    9'd347: begin
      dout <= mem_space[347];
    end
    9'd348: begin
      dout <= mem_space[348];
    end
    9'd349: begin
      dout <= mem_space[349];
    end
    9'd350: begin
      dout <= mem_space[350];
    end
    9'd351: begin
      dout <= mem_space[351];
    end
    9'd352: begin
      dout <= mem_space[352];
    end
    9'd353: begin
      dout <= mem_space[353];
    end
    9'd354: begin
      dout <= mem_space[354];
    end
    9'd355: begin
      dout <= mem_space[355];
    end
    9'd356: begin
      dout <= mem_space[356];
    end
    9'd357: begin
      dout <= mem_space[357];
    end
    9'd358: begin
      dout <= mem_space[358];
    end
    9'd359: begin
      dout <= mem_space[359];
    end
    9'd360: begin
      dout <= mem_space[360];
    end
    9'd361: begin
      dout <= mem_space[361];
    end
    9'd362: begin
      dout <= mem_space[362];
    end
    9'd363: begin
      dout <= mem_space[363];
    end
    9'd364: begin
      dout <= mem_space[364];
    end
    9'd365: begin
      dout <= mem_space[365];
    end
    9'd366: begin
      dout <= mem_space[366];
    end
    9'd367: begin
      dout <= mem_space[367];
    end
    9'd368: begin
      dout <= mem_space[368];
    end
    9'd369: begin
      dout <= mem_space[369];
    end
    9'd370: begin
      dout <= mem_space[370];
    end
    9'd371: begin
      dout <= mem_space[371];
    end
    9'd372: begin
      dout <= mem_space[372];
    end
    9'd373: begin
      dout <= mem_space[373];
    end
    9'd374: begin
      dout <= mem_space[374];
    end
    9'd375: begin
      dout <= mem_space[375];
    end
    9'd376: begin
      dout <= mem_space[376];
    end
    9'd377: begin
      dout <= mem_space[377];
    end
    9'd378: begin
      dout <= mem_space[378];
    end
    9'd379: begin
      dout <= mem_space[379];
    end
    9'd380: begin
      dout <= mem_space[380];
    end
    9'd381: begin
      dout <= mem_space[381];
    end
    9'd382: begin
      dout <= mem_space[382];
    end
    9'd383: begin
      dout <= mem_space[383];
    end
    9'd384: begin
      dout <= mem_space[384];
    end
    9'd385: begin
      dout <= mem_space[385];
    end
    9'd386: begin
      dout <= mem_space[386];
    end
    9'd387: begin
      dout <= mem_space[387];
    end
    9'd388: begin
      dout <= mem_space[388];
    end
    9'd389: begin
      dout <= mem_space[389];
    end
    9'd390: begin
      dout <= mem_space[390];
    end
    9'd391: begin
      dout <= mem_space[391];
    end
    9'd392: begin
      dout <= mem_space[392];
    end
    9'd393: begin
      dout <= mem_space[393];
    end
    9'd394: begin
      dout <= mem_space[394];
    end
    9'd395: begin
      dout <= mem_space[395];
    end
    9'd396: begin
      dout <= mem_space[396];
    end
    9'd397: begin
      dout <= mem_space[397];
    end
    9'd398: begin
      dout <= mem_space[398];
    end
    9'd399: begin
      dout <= mem_space[399];
    end
    9'd400: begin
      dout <= mem_space[400];
    end
    9'd401: begin
      dout <= mem_space[401];
    end
    9'd402: begin
      dout <= mem_space[402];
    end
    9'd403: begin
      dout <= mem_space[403];
    end
    9'd404: begin
      dout <= mem_space[404];
    end
    9'd405: begin
      dout <= mem_space[405];
    end
    9'd406: begin
      dout <= mem_space[406];
    end
    9'd407: begin
      dout <= mem_space[407];
    end
    9'd408: begin
      dout <= mem_space[408];
    end
    9'd409: begin
      dout <= mem_space[409];
    end
    9'd410: begin
      dout <= mem_space[410];
    end
    9'd411: begin
      dout <= mem_space[411];
    end
    9'd412: begin
      dout <= mem_space[412];
    end
    9'd413: begin
      dout <= mem_space[413];
    end
    9'd414: begin
      dout <= mem_space[414];
    end
    9'd415: begin
      dout <= mem_space[415];
    end
    9'd416: begin
      dout <= mem_space[416];
    end
    9'd417: begin
      dout <= mem_space[417];
    end
    9'd418: begin
      dout <= mem_space[418];
    end
    9'd419: begin
      dout <= mem_space[419];
    end
    9'd420: begin
      dout <= mem_space[420];
    end
    9'd421: begin
      dout <= mem_space[421];
    end
    9'd422: begin
      dout <= mem_space[422];
    end
    9'd423: begin
      dout <= mem_space[423];
    end
    9'd424: begin
      dout <= mem_space[424];
    end
    9'd425: begin
      dout <= mem_space[425];
    end
    9'd426: begin
      dout <= mem_space[426];
    end
    9'd427: begin
      dout <= mem_space[427];
    end
    9'd428: begin
      dout <= mem_space[428];
    end
    9'd429: begin
      dout <= mem_space[429];
    end
    9'd430: begin
      dout <= mem_space[430];
    end
    9'd431: begin
      dout <= mem_space[431];
    end
    9'd432: begin
      dout <= mem_space[432];
    end
    9'd433: begin
      dout <= mem_space[433];
    end
    9'd434: begin
      dout <= mem_space[434];
    end
    9'd435: begin
      dout <= mem_space[435];
    end
    9'd436: begin
      dout <= mem_space[436];
    end
    9'd437: begin
      dout <= mem_space[437];
    end
    9'd438: begin
      dout <= mem_space[438];
    end
    9'd439: begin
      dout <= mem_space[439];
    end
    9'd440: begin
      dout <= mem_space[440];
    end
    9'd441: begin
      dout <= mem_space[441];
    end
    9'd442: begin
      dout <= mem_space[442];
    end
    9'd443: begin
      dout <= mem_space[443];
    end
    9'd444: begin
      dout <= mem_space[444];
    end
    9'd445: begin
      dout <= mem_space[445];
    end
    9'd446: begin
      dout <= mem_space[446];
    end
    9'd447: begin
      dout <= mem_space[447];
    end
    9'd448: begin
      dout <= mem_space[448];
    end
    9'd449: begin
      dout <= mem_space[449];
    end
    9'd450: begin
      dout <= mem_space[450];
    end
    9'd451: begin
      dout <= mem_space[451];
    end
    9'd452: begin
      dout <= mem_space[452];
    end
    9'd453: begin
      dout <= mem_space[453];
    end
    9'd454: begin
      dout <= mem_space[454];
    end
    9'd455: begin
      dout <= mem_space[455];
    end
    9'd456: begin
      dout <= mem_space[456];
    end
    9'd457: begin
      dout <= mem_space[457];
    end
    9'd458: begin
      dout <= mem_space[458];
    end
    9'd459: begin
      dout <= mem_space[459];
    end
    9'd460: begin
      dout <= mem_space[460];
    end
    9'd461: begin
      dout <= mem_space[461];
    end
    9'd462: begin
      dout <= mem_space[462];
    end
    9'd463: begin
      dout <= mem_space[463];
    end
    9'd464: begin
      dout <= mem_space[464];
    end
    9'd465: begin
      dout <= mem_space[465];
    end
    9'd466: begin
      dout <= mem_space[466];
    end
    9'd467: begin
      dout <= mem_space[467];
    end
    9'd468: begin
      dout <= mem_space[468];
    end
    9'd469: begin
      dout <= mem_space[469];
    end
    9'd470: begin
      dout <= mem_space[470];
    end
    9'd471: begin
      dout <= mem_space[471];
    end
    9'd472: begin
      dout <= mem_space[472];
    end
    9'd473: begin
      dout <= mem_space[473];
    end
    9'd474: begin
      dout <= mem_space[474];
    end
    9'd475: begin
      dout <= mem_space[475];
    end
    9'd476: begin
      dout <= mem_space[476];
    end
    9'd477: begin
      dout <= mem_space[477];
    end
    9'd478: begin
      dout <= mem_space[478];
    end
    9'd479: begin
      dout <= mem_space[479];
    end
    9'd480: begin
      dout <= mem_space[480];
    end
    9'd481: begin
      dout <= mem_space[481];
    end
    9'd482: begin
      dout <= mem_space[482];
    end
    9'd483: begin
      dout <= mem_space[483];
    end
    9'd484: begin
      dout <= mem_space[484];
    end
    9'd485: begin
      dout <= mem_space[485];
    end
    9'd486: begin
      dout <= mem_space[486];
    end
    9'd487: begin
      dout <= mem_space[487];
    end
    9'd488: begin
      dout <= mem_space[488];
    end
    9'd489: begin
      dout <= mem_space[489];
    end
    9'd490: begin
      dout <= mem_space[490];
    end
    9'd491: begin
      dout <= mem_space[491];
    end
    9'd492: begin
      dout <= mem_space[492];
    end
    9'd493: begin
      dout <= mem_space[493];
    end
    9'd494: begin
      dout <= mem_space[494];
    end
    9'd495: begin
      dout <= mem_space[495];
    end
    9'd496: begin
      dout <= mem_space[496];
    end
    9'd497: begin
      dout <= mem_space[497];
    end
    9'd498: begin
      dout <= mem_space[498];
    end
    9'd499: begin
      dout <= mem_space[499];
    end
    9'd500: begin
      dout <= mem_space[500];
    end
    9'd501: begin
      dout <= mem_space[501];
    end
    9'd502: begin
      dout <= mem_space[502];
    end
    9'd503: begin
      dout <= mem_space[503];
    end
    9'd504: begin
      dout <= mem_space[504];
    end
    9'd505: begin
      dout <= mem_space[505];
    end
    9'd506: begin
      dout <= mem_space[506];
    end
    9'd507: begin
      dout <= mem_space[507];
    end
    9'd508: begin
      dout <= mem_space[508];
    end
    9'd509: begin
      dout <= mem_space[509];
    end
    9'd510: begin
      dout <= mem_space[510];
    end
    9'd511: begin
      dout <= mem_space[511];
    end
  endcase
end

always_ff@(posedge clk) begin
  case( raddr )
    9'd0: begin
     mem_space[0] <= din;
    end
    9'd1: begin
     mem_space[1] <= din;
    end
    9'd2: begin
     mem_space[2] <= din;
    end
    9'd3: begin
     mem_space[3] <= din;
    end
    9'd4: begin
     mem_space[4] <= din;
    end
    9'd5: begin
     mem_space[5] <= din;
    end
    9'd6: begin
     mem_space[6] <= din;
    end
    9'd7: begin
     mem_space[7] <= din;
    end
    9'd8: begin
     mem_space[8] <= din;
    end
    9'd9: begin
     mem_space[9] <= din;
    end
    9'd10: begin
     mem_space[10] <= din;
    end
    9'd11: begin
     mem_space[11] <= din;
    end
    9'd12: begin
     mem_space[12] <= din;
    end
    9'd13: begin
     mem_space[13] <= din;
    end
    9'd14: begin
     mem_space[14] <= din;
    end
    9'd15: begin
     mem_space[15] <= din;
    end
    9'd16: begin
     mem_space[16] <= din;
    end
    9'd17: begin
     mem_space[17] <= din;
    end
    9'd18: begin
     mem_space[18] <= din;
    end
    9'd19: begin
     mem_space[19] <= din;
    end
    9'd20: begin
     mem_space[20] <= din;
    end
    9'd21: begin
     mem_space[21] <= din;
    end
    9'd22: begin
     mem_space[22] <= din;
    end
    9'd23: begin
     mem_space[23] <= din;
    end
    9'd24: begin
     mem_space[24] <= din;
    end
    9'd25: begin
     mem_space[25] <= din;
    end
    9'd26: begin
     mem_space[26] <= din;
    end
    9'd27: begin
     mem_space[27] <= din;
    end
    9'd28: begin
     mem_space[28] <= din;
    end
    9'd29: begin
     mem_space[29] <= din;
    end
    9'd30: begin
     mem_space[30] <= din;
    end
    9'd31: begin
     mem_space[31] <= din;
    end
    9'd32: begin
     mem_space[32] <= din;
    end
    9'd33: begin
     mem_space[33] <= din;
    end
    9'd34: begin
     mem_space[34] <= din;
    end
    9'd35: begin
     mem_space[35] <= din;
    end
    9'd36: begin
     mem_space[36] <= din;
    end
    9'd37: begin
     mem_space[37] <= din;
    end
    9'd38: begin
     mem_space[38] <= din;
    end
    9'd39: begin
     mem_space[39] <= din;
    end
    9'd40: begin
     mem_space[40] <= din;
    end
    9'd41: begin
     mem_space[41] <= din;
    end
    9'd42: begin
     mem_space[42] <= din;
    end
    9'd43: begin
     mem_space[43] <= din;
    end
    9'd44: begin
     mem_space[44] <= din;
    end
    9'd45: begin
     mem_space[45] <= din;
    end
    9'd46: begin
     mem_space[46] <= din;
    end
    9'd47: begin
     mem_space[47] <= din;
    end
    9'd48: begin
     mem_space[48] <= din;
    end
    9'd49: begin
     mem_space[49] <= din;
    end
    9'd50: begin
     mem_space[50] <= din;
    end
    9'd51: begin
     mem_space[51] <= din;
    end
    9'd52: begin
     mem_space[52] <= din;
    end
    9'd53: begin
     mem_space[53] <= din;
    end
    9'd54: begin
     mem_space[54] <= din;
    end
    9'd55: begin
     mem_space[55] <= din;
    end
    9'd56: begin
     mem_space[56] <= din;
    end
    9'd57: begin
     mem_space[57] <= din;
    end
    9'd58: begin
     mem_space[58] <= din;
    end
    9'd59: begin
     mem_space[59] <= din;
    end
    9'd60: begin
     mem_space[60] <= din;
    end
    9'd61: begin
     mem_space[61] <= din;
    end
    9'd62: begin
     mem_space[62] <= din;
    end
    9'd63: begin
     mem_space[63] <= din;
    end
    9'd64: begin
     mem_space[64] <= din;
    end
    9'd65: begin
     mem_space[65] <= din;
    end
    9'd66: begin
     mem_space[66] <= din;
    end
    9'd67: begin
     mem_space[67] <= din;
    end
    9'd68: begin
     mem_space[68] <= din;
    end
    9'd69: begin
     mem_space[69] <= din;
    end
    9'd70: begin
     mem_space[70] <= din;
    end
    9'd71: begin
     mem_space[71] <= din;
    end
    9'd72: begin
     mem_space[72] <= din;
    end
    9'd73: begin
     mem_space[73] <= din;
    end
    9'd74: begin
     mem_space[74] <= din;
    end
    9'd75: begin
     mem_space[75] <= din;
    end
    9'd76: begin
     mem_space[76] <= din;
    end
    9'd77: begin
     mem_space[77] <= din;
    end
    9'd78: begin
     mem_space[78] <= din;
    end
    9'd79: begin
     mem_space[79] <= din;
    end
    9'd80: begin
     mem_space[80] <= din;
    end
    9'd81: begin
     mem_space[81] <= din;
    end
    9'd82: begin
     mem_space[82] <= din;
    end
    9'd83: begin
     mem_space[83] <= din;
    end
    9'd84: begin
     mem_space[84] <= din;
    end
    9'd85: begin
     mem_space[85] <= din;
    end
    9'd86: begin
     mem_space[86] <= din;
    end
    9'd87: begin
     mem_space[87] <= din;
    end
    9'd88: begin
     mem_space[88] <= din;
    end
    9'd89: begin
     mem_space[89] <= din;
    end
    9'd90: begin
     mem_space[90] <= din;
    end
    9'd91: begin
     mem_space[91] <= din;
    end
    9'd92: begin
     mem_space[92] <= din;
    end
    9'd93: begin
     mem_space[93] <= din;
    end
    9'd94: begin
     mem_space[94] <= din;
    end
    9'd95: begin
     mem_space[95] <= din;
    end
    9'd96: begin
     mem_space[96] <= din;
    end
    9'd97: begin
     mem_space[97] <= din;
    end
    9'd98: begin
     mem_space[98] <= din;
    end
    9'd99: begin
     mem_space[99] <= din;
    end
    9'd100: begin
     mem_space[100] <= din;
    end
    9'd101: begin
     mem_space[101] <= din;
    end
    9'd102: begin
     mem_space[102] <= din;
    end
    9'd103: begin
     mem_space[103] <= din;
    end
    9'd104: begin
     mem_space[104] <= din;
    end
    9'd105: begin
     mem_space[105] <= din;
    end
    9'd106: begin
     mem_space[106] <= din;
    end
    9'd107: begin
     mem_space[107] <= din;
    end
    9'd108: begin
     mem_space[108] <= din;
    end
    9'd109: begin
     mem_space[109] <= din;
    end
    9'd110: begin
     mem_space[110] <= din;
    end
    9'd111: begin
     mem_space[111] <= din;
    end
    9'd112: begin
     mem_space[112] <= din;
    end
    9'd113: begin
     mem_space[113] <= din;
    end
    9'd114: begin
     mem_space[114] <= din;
    end
    9'd115: begin
     mem_space[115] <= din;
    end
    9'd116: begin
     mem_space[116] <= din;
    end
    9'd117: begin
     mem_space[117] <= din;
    end
    9'd118: begin
     mem_space[118] <= din;
    end
    9'd119: begin
     mem_space[119] <= din;
    end
    9'd120: begin
     mem_space[120] <= din;
    end
    9'd121: begin
     mem_space[121] <= din;
    end
    9'd122: begin
     mem_space[122] <= din;
    end
    9'd123: begin
     mem_space[123] <= din;
    end
    9'd124: begin
     mem_space[124] <= din;
    end
    9'd125: begin
     mem_space[125] <= din;
    end
    9'd126: begin
     mem_space[126] <= din;
    end
    9'd127: begin
     mem_space[127] <= din;
    end
    9'd128: begin
     mem_space[128] <= din;
    end
    9'd129: begin
     mem_space[129] <= din;
    end
    9'd130: begin
     mem_space[130] <= din;
    end
    9'd131: begin
     mem_space[131] <= din;
    end
    9'd132: begin
     mem_space[132] <= din;
    end
    9'd133: begin
     mem_space[133] <= din;
    end
    9'd134: begin
     mem_space[134] <= din;
    end
    9'd135: begin
     mem_space[135] <= din;
    end
    9'd136: begin
     mem_space[136] <= din;
    end
    9'd137: begin
     mem_space[137] <= din;
    end
    9'd138: begin
     mem_space[138] <= din;
    end
    9'd139: begin
     mem_space[139] <= din;
    end
    9'd140: begin
     mem_space[140] <= din;
    end
    9'd141: begin
     mem_space[141] <= din;
    end
    9'd142: begin
     mem_space[142] <= din;
    end
    9'd143: begin
     mem_space[143] <= din;
    end
    9'd144: begin
     mem_space[144] <= din;
    end
    9'd145: begin
     mem_space[145] <= din;
    end
    9'd146: begin
     mem_space[146] <= din;
    end
    9'd147: begin
     mem_space[147] <= din;
    end
    9'd148: begin
     mem_space[148] <= din;
    end
    9'd149: begin
     mem_space[149] <= din;
    end
    9'd150: begin
     mem_space[150] <= din;
    end
    9'd151: begin
     mem_space[151] <= din;
    end
    9'd152: begin
     mem_space[152] <= din;
    end
    9'd153: begin
     mem_space[153] <= din;
    end
    9'd154: begin
     mem_space[154] <= din;
    end
    9'd155: begin
     mem_space[155] <= din;
    end
    9'd156: begin
     mem_space[156] <= din;
    end
    9'd157: begin
     mem_space[157] <= din;
    end
    9'd158: begin
     mem_space[158] <= din;
    end
    9'd159: begin
     mem_space[159] <= din;
    end
    9'd160: begin
     mem_space[160] <= din;
    end
    9'd161: begin
     mem_space[161] <= din;
    end
    9'd162: begin
     mem_space[162] <= din;
    end
    9'd163: begin
     mem_space[163] <= din;
    end
    9'd164: begin
     mem_space[164] <= din;
    end
    9'd165: begin
     mem_space[165] <= din;
    end
    9'd166: begin
     mem_space[166] <= din;
    end
    9'd167: begin
     mem_space[167] <= din;
    end
    9'd168: begin
     mem_space[168] <= din;
    end
    9'd169: begin
     mem_space[169] <= din;
    end
    9'd170: begin
     mem_space[170] <= din;
    end
    9'd171: begin
     mem_space[171] <= din;
    end
    9'd172: begin
     mem_space[172] <= din;
    end
    9'd173: begin
     mem_space[173] <= din;
    end
    9'd174: begin
     mem_space[174] <= din;
    end
    9'd175: begin
     mem_space[175] <= din;
    end
    9'd176: begin
     mem_space[176] <= din;
    end
    9'd177: begin
     mem_space[177] <= din;
    end
    9'd178: begin
     mem_space[178] <= din;
    end
    9'd179: begin
     mem_space[179] <= din;
    end
    9'd180: begin
     mem_space[180] <= din;
    end
    9'd181: begin
     mem_space[181] <= din;
    end
    9'd182: begin
     mem_space[182] <= din;
    end
    9'd183: begin
     mem_space[183] <= din;
    end
    9'd184: begin
     mem_space[184] <= din;
    end
    9'd185: begin
     mem_space[185] <= din;
    end
    9'd186: begin
     mem_space[186] <= din;
    end
    9'd187: begin
     mem_space[187] <= din;
    end
    9'd188: begin
     mem_space[188] <= din;
    end
    9'd189: begin
     mem_space[189] <= din;
    end
    9'd190: begin
     mem_space[190] <= din;
    end
    9'd191: begin
     mem_space[191] <= din;
    end
    9'd192: begin
     mem_space[192] <= din;
    end
    9'd193: begin
     mem_space[193] <= din;
    end
    9'd194: begin
     mem_space[194] <= din;
    end
    9'd195: begin
     mem_space[195] <= din;
    end
    9'd196: begin
     mem_space[196] <= din;
    end
    9'd197: begin
     mem_space[197] <= din;
    end
    9'd198: begin
     mem_space[198] <= din;
    end
    9'd199: begin
     mem_space[199] <= din;
    end
    9'd200: begin
     mem_space[200] <= din;
    end
    9'd201: begin
     mem_space[201] <= din;
    end
    9'd202: begin
     mem_space[202] <= din;
    end
    9'd203: begin
     mem_space[203] <= din;
    end
    9'd204: begin
     mem_space[204] <= din;
    end
    9'd205: begin
     mem_space[205] <= din;
    end
    9'd206: begin
     mem_space[206] <= din;
    end
    9'd207: begin
     mem_space[207] <= din;
    end
    9'd208: begin
     mem_space[208] <= din;
    end
    9'd209: begin
     mem_space[209] <= din;
    end
    9'd210: begin
     mem_space[210] <= din;
    end
    9'd211: begin
     mem_space[211] <= din;
    end
    9'd212: begin
     mem_space[212] <= din;
    end
    9'd213: begin
     mem_space[213] <= din;
    end
    9'd214: begin
     mem_space[214] <= din;
    end
    9'd215: begin
     mem_space[215] <= din;
    end
    9'd216: begin
     mem_space[216] <= din;
    end
    9'd217: begin
     mem_space[217] <= din;
    end
    9'd218: begin
     mem_space[218] <= din;
    end
    9'd219: begin
     mem_space[219] <= din;
    end
    9'd220: begin
     mem_space[220] <= din;
    end
    9'd221: begin
     mem_space[221] <= din;
    end
    9'd222: begin
     mem_space[222] <= din;
    end
    9'd223: begin
     mem_space[223] <= din;
    end
    9'd224: begin
     mem_space[224] <= din;
    end
    9'd225: begin
     mem_space[225] <= din;
    end
    9'd226: begin
     mem_space[226] <= din;
    end
    9'd227: begin
     mem_space[227] <= din;
    end
    9'd228: begin
     mem_space[228] <= din;
    end
    9'd229: begin
     mem_space[229] <= din;
    end
    9'd230: begin
     mem_space[230] <= din;
    end
    9'd231: begin
     mem_space[231] <= din;
    end
    9'd232: begin
     mem_space[232] <= din;
    end
    9'd233: begin
     mem_space[233] <= din;
    end
    9'd234: begin
     mem_space[234] <= din;
    end
    9'd235: begin
     mem_space[235] <= din;
    end
    9'd236: begin
     mem_space[236] <= din;
    end
    9'd237: begin
     mem_space[237] <= din;
    end
    9'd238: begin
     mem_space[238] <= din;
    end
    9'd239: begin
     mem_space[239] <= din;
    end
    9'd240: begin
     mem_space[240] <= din;
    end
    9'd241: begin
     mem_space[241] <= din;
    end
    9'd242: begin
     mem_space[242] <= din;
    end
    9'd243: begin
     mem_space[243] <= din;
    end
    9'd244: begin
     mem_space[244] <= din;
    end
    9'd245: begin
     mem_space[245] <= din;
    end
    9'd246: begin
     mem_space[246] <= din;
    end
    9'd247: begin
     mem_space[247] <= din;
    end
    9'd248: begin
     mem_space[248] <= din;
    end
    9'd249: begin
     mem_space[249] <= din;
    end
    9'd250: begin
     mem_space[250] <= din;
    end
    9'd251: begin
     mem_space[251] <= din;
    end
    9'd252: begin
     mem_space[252] <= din;
    end
    9'd253: begin
     mem_space[253] <= din;
    end
    9'd254: begin
     mem_space[254] <= din;
    end
    9'd255: begin
     mem_space[255] <= din;
    end
    9'd256: begin
     mem_space[256] <= din;
    end
    9'd257: begin
     mem_space[257] <= din;
    end
    9'd258: begin
     mem_space[258] <= din;
    end
    9'd259: begin
     mem_space[259] <= din;
    end
    9'd260: begin
     mem_space[260] <= din;
    end
    9'd261: begin
     mem_space[261] <= din;
    end
    9'd262: begin
     mem_space[262] <= din;
    end
    9'd263: begin
     mem_space[263] <= din;
    end
    9'd264: begin
     mem_space[264] <= din;
    end
    9'd265: begin
     mem_space[265] <= din;
    end
    9'd266: begin
     mem_space[266] <= din;
    end
    9'd267: begin
     mem_space[267] <= din;
    end
    9'd268: begin
     mem_space[268] <= din;
    end
    9'd269: begin
     mem_space[269] <= din;
    end
    9'd270: begin
     mem_space[270] <= din;
    end
    9'd271: begin
     mem_space[271] <= din;
    end
    9'd272: begin
     mem_space[272] <= din;
    end
    9'd273: begin
     mem_space[273] <= din;
    end
    9'd274: begin
     mem_space[274] <= din;
    end
    9'd275: begin
     mem_space[275] <= din;
    end
    9'd276: begin
     mem_space[276] <= din;
    end
    9'd277: begin
     mem_space[277] <= din;
    end
    9'd278: begin
     mem_space[278] <= din;
    end
    9'd279: begin
     mem_space[279] <= din;
    end
    9'd280: begin
     mem_space[280] <= din;
    end
    9'd281: begin
     mem_space[281] <= din;
    end
    9'd282: begin
     mem_space[282] <= din;
    end
    9'd283: begin
     mem_space[283] <= din;
    end
    9'd284: begin
     mem_space[284] <= din;
    end
    9'd285: begin
     mem_space[285] <= din;
    end
    9'd286: begin
     mem_space[286] <= din;
    end
    9'd287: begin
     mem_space[287] <= din;
    end
    9'd288: begin
     mem_space[288] <= din;
    end
    9'd289: begin
     mem_space[289] <= din;
    end
    9'd290: begin
     mem_space[290] <= din;
    end
    9'd291: begin
     mem_space[291] <= din;
    end
    9'd292: begin
     mem_space[292] <= din;
    end
    9'd293: begin
     mem_space[293] <= din;
    end
    9'd294: begin
     mem_space[294] <= din;
    end
    9'd295: begin
     mem_space[295] <= din;
    end
    9'd296: begin
     mem_space[296] <= din;
    end
    9'd297: begin
     mem_space[297] <= din;
    end
    9'd298: begin
     mem_space[298] <= din;
    end
    9'd299: begin
     mem_space[299] <= din;
    end
    9'd300: begin
     mem_space[300] <= din;
    end
    9'd301: begin
     mem_space[301] <= din;
    end
    9'd302: begin
     mem_space[302] <= din;
    end
    9'd303: begin
     mem_space[303] <= din;
    end
    9'd304: begin
     mem_space[304] <= din;
    end
    9'd305: begin
     mem_space[305] <= din;
    end
    9'd306: begin
     mem_space[306] <= din;
    end
    9'd307: begin
     mem_space[307] <= din;
    end
    9'd308: begin
     mem_space[308] <= din;
    end
    9'd309: begin
     mem_space[309] <= din;
    end
    9'd310: begin
     mem_space[310] <= din;
    end
    9'd311: begin
     mem_space[311] <= din;
    end
    9'd312: begin
     mem_space[312] <= din;
    end
    9'd313: begin
     mem_space[313] <= din;
    end
    9'd314: begin
     mem_space[314] <= din;
    end
    9'd315: begin
     mem_space[315] <= din;
    end
    9'd316: begin
     mem_space[316] <= din;
    end
    9'd317: begin
     mem_space[317] <= din;
    end
    9'd318: begin
     mem_space[318] <= din;
    end
    9'd319: begin
     mem_space[319] <= din;
    end
    9'd320: begin
     mem_space[320] <= din;
    end
    9'd321: begin
     mem_space[321] <= din;
    end
    9'd322: begin
     mem_space[322] <= din;
    end
    9'd323: begin
     mem_space[323] <= din;
    end
    9'd324: begin
     mem_space[324] <= din;
    end
    9'd325: begin
     mem_space[325] <= din;
    end
    9'd326: begin
     mem_space[326] <= din;
    end
    9'd327: begin
     mem_space[327] <= din;
    end
    9'd328: begin
     mem_space[328] <= din;
    end
    9'd329: begin
     mem_space[329] <= din;
    end
    9'd330: begin
     mem_space[330] <= din;
    end
    9'd331: begin
     mem_space[331] <= din;
    end
    9'd332: begin
     mem_space[332] <= din;
    end
    9'd333: begin
     mem_space[333] <= din;
    end
    9'd334: begin
     mem_space[334] <= din;
    end
    9'd335: begin
     mem_space[335] <= din;
    end
    9'd336: begin
     mem_space[336] <= din;
    end
    9'd337: begin
     mem_space[337] <= din;
    end
    9'd338: begin
     mem_space[338] <= din;
    end
    9'd339: begin
     mem_space[339] <= din;
    end
    9'd340: begin
     mem_space[340] <= din;
    end
    9'd341: begin
     mem_space[341] <= din;
    end
    9'd342: begin
     mem_space[342] <= din;
    end
    9'd343: begin
     mem_space[343] <= din;
    end
    9'd344: begin
     mem_space[344] <= din;
    end
    9'd345: begin
     mem_space[345] <= din;
    end
    9'd346: begin
     mem_space[346] <= din;
    end
    9'd347: begin
     mem_space[347] <= din;
    end
    9'd348: begin
     mem_space[348] <= din;
    end
    9'd349: begin
     mem_space[349] <= din;
    end
    9'd350: begin
     mem_space[350] <= din;
    end
    9'd351: begin
     mem_space[351] <= din;
    end
    9'd352: begin
     mem_space[352] <= din;
    end
    9'd353: begin
     mem_space[353] <= din;
    end
    9'd354: begin
     mem_space[354] <= din;
    end
    9'd355: begin
     mem_space[355] <= din;
    end
    9'd356: begin
     mem_space[356] <= din;
    end
    9'd357: begin
     mem_space[357] <= din;
    end
    9'd358: begin
     mem_space[358] <= din;
    end
    9'd359: begin
     mem_space[359] <= din;
    end
    9'd360: begin
     mem_space[360] <= din;
    end
    9'd361: begin
     mem_space[361] <= din;
    end
    9'd362: begin
     mem_space[362] <= din;
    end
    9'd363: begin
     mem_space[363] <= din;
    end
    9'd364: begin
     mem_space[364] <= din;
    end
    9'd365: begin
     mem_space[365] <= din;
    end
    9'd366: begin
     mem_space[366] <= din;
    end
    9'd367: begin
     mem_space[367] <= din;
    end
    9'd368: begin
     mem_space[368] <= din;
    end
    9'd369: begin
     mem_space[369] <= din;
    end
    9'd370: begin
     mem_space[370] <= din;
    end
    9'd371: begin
     mem_space[371] <= din;
    end
    9'd372: begin
     mem_space[372] <= din;
    end
    9'd373: begin
     mem_space[373] <= din;
    end
    9'd374: begin
     mem_space[374] <= din;
    end
    9'd375: begin
     mem_space[375] <= din;
    end
    9'd376: begin
     mem_space[376] <= din;
    end
    9'd377: begin
     mem_space[377] <= din;
    end
    9'd378: begin
     mem_space[378] <= din;
    end
    9'd379: begin
     mem_space[379] <= din;
    end
    9'd380: begin
     mem_space[380] <= din;
    end
    9'd381: begin
     mem_space[381] <= din;
    end
    9'd382: begin
     mem_space[382] <= din;
    end
    9'd383: begin
     mem_space[383] <= din;
    end
    9'd384: begin
     mem_space[384] <= din;
    end
    9'd385: begin
     mem_space[385] <= din;
    end
    9'd386: begin
     mem_space[386] <= din;
    end
    9'd387: begin
     mem_space[387] <= din;
    end
    9'd388: begin
     mem_space[388] <= din;
    end
    9'd389: begin
     mem_space[389] <= din;
    end
    9'd390: begin
     mem_space[390] <= din;
    end
    9'd391: begin
     mem_space[391] <= din;
    end
    9'd392: begin
     mem_space[392] <= din;
    end
    9'd393: begin
     mem_space[393] <= din;
    end
    9'd394: begin
     mem_space[394] <= din;
    end
    9'd395: begin
     mem_space[395] <= din;
    end
    9'd396: begin
     mem_space[396] <= din;
    end
    9'd397: begin
     mem_space[397] <= din;
    end
    9'd398: begin
     mem_space[398] <= din;
    end
    9'd399: begin
     mem_space[399] <= din;
    end
    9'd400: begin
     mem_space[400] <= din;
    end
    9'd401: begin
     mem_space[401] <= din;
    end
    9'd402: begin
     mem_space[402] <= din;
    end
    9'd403: begin
     mem_space[403] <= din;
    end
    9'd404: begin
     mem_space[404] <= din;
    end
    9'd405: begin
     mem_space[405] <= din;
    end
    9'd406: begin
     mem_space[406] <= din;
    end
    9'd407: begin
     mem_space[407] <= din;
    end
    9'd408: begin
     mem_space[408] <= din;
    end
    9'd409: begin
     mem_space[409] <= din;
    end
    9'd410: begin
     mem_space[410] <= din;
    end
    9'd411: begin
     mem_space[411] <= din;
    end
    9'd412: begin
     mem_space[412] <= din;
    end
    9'd413: begin
     mem_space[413] <= din;
    end
    9'd414: begin
     mem_space[414] <= din;
    end
    9'd415: begin
     mem_space[415] <= din;
    end
    9'd416: begin
     mem_space[416] <= din;
    end
    9'd417: begin
     mem_space[417] <= din;
    end
    9'd418: begin
     mem_space[418] <= din;
    end
    9'd419: begin
     mem_space[419] <= din;
    end
    9'd420: begin
     mem_space[420] <= din;
    end
    9'd421: begin
     mem_space[421] <= din;
    end
    9'd422: begin
     mem_space[422] <= din;
    end
    9'd423: begin
     mem_space[423] <= din;
    end
    9'd424: begin
     mem_space[424] <= din;
    end
    9'd425: begin
     mem_space[425] <= din;
    end
    9'd426: begin
     mem_space[426] <= din;
    end
    9'd427: begin
     mem_space[427] <= din;
    end
    9'd428: begin
     mem_space[428] <= din;
    end
    9'd429: begin
     mem_space[429] <= din;
    end
    9'd430: begin
     mem_space[430] <= din;
    end
    9'd431: begin
     mem_space[431] <= din;
    end
    9'd432: begin
     mem_space[432] <= din;
    end
    9'd433: begin
     mem_space[433] <= din;
    end
    9'd434: begin
     mem_space[434] <= din;
    end
    9'd435: begin
     mem_space[435] <= din;
    end
    9'd436: begin
     mem_space[436] <= din;
    end
    9'd437: begin
     mem_space[437] <= din;
    end
    9'd438: begin
     mem_space[438] <= din;
    end
    9'd439: begin
     mem_space[439] <= din;
    end
    9'd440: begin
     mem_space[440] <= din;
    end
    9'd441: begin
     mem_space[441] <= din;
    end
    9'd442: begin
     mem_space[442] <= din;
    end
    9'd443: begin
     mem_space[443] <= din;
    end
    9'd444: begin
     mem_space[444] <= din;
    end
    9'd445: begin
     mem_space[445] <= din;
    end
    9'd446: begin
     mem_space[446] <= din;
    end
    9'd447: begin
     mem_space[447] <= din;
    end
    9'd448: begin
     mem_space[448] <= din;
    end
    9'd449: begin
     mem_space[449] <= din;
    end
    9'd450: begin
     mem_space[450] <= din;
    end
    9'd451: begin
     mem_space[451] <= din;
    end
    9'd452: begin
     mem_space[452] <= din;
    end
    9'd453: begin
     mem_space[453] <= din;
    end
    9'd454: begin
     mem_space[454] <= din;
    end
    9'd455: begin
     mem_space[455] <= din;
    end
    9'd456: begin
     mem_space[456] <= din;
    end
    9'd457: begin
     mem_space[457] <= din;
    end
    9'd458: begin
     mem_space[458] <= din;
    end
    9'd459: begin
     mem_space[459] <= din;
    end
    9'd460: begin
     mem_space[460] <= din;
    end
    9'd461: begin
     mem_space[461] <= din;
    end
    9'd462: begin
     mem_space[462] <= din;
    end
    9'd463: begin
     mem_space[463] <= din;
    end
    9'd464: begin
     mem_space[464] <= din;
    end
    9'd465: begin
     mem_space[465] <= din;
    end
    9'd466: begin
     mem_space[466] <= din;
    end
    9'd467: begin
     mem_space[467] <= din;
    end
    9'd468: begin
     mem_space[468] <= din;
    end
    9'd469: begin
     mem_space[469] <= din;
    end
    9'd470: begin
     mem_space[470] <= din;
    end
    9'd471: begin
     mem_space[471] <= din;
    end
    9'd472: begin
     mem_space[472] <= din;
    end
    9'd473: begin
     mem_space[473] <= din;
    end
    9'd474: begin
     mem_space[474] <= din;
    end
    9'd475: begin
     mem_space[475] <= din;
    end
    9'd476: begin
     mem_space[476] <= din;
    end
    9'd477: begin
     mem_space[477] <= din;
    end
    9'd478: begin
     mem_space[478] <= din;
    end
    9'd479: begin
     mem_space[479] <= din;
    end
    9'd480: begin
     mem_space[480] <= din;
    end
    9'd481: begin
     mem_space[481] <= din;
    end
    9'd482: begin
     mem_space[482] <= din;
    end
    9'd483: begin
     mem_space[483] <= din;
    end
    9'd484: begin
     mem_space[484] <= din;
    end
    9'd485: begin
     mem_space[485] <= din;
    end
    9'd486: begin
     mem_space[486] <= din;
    end
    9'd487: begin
     mem_space[487] <= din;
    end
    9'd488: begin
     mem_space[488] <= din;
    end
    9'd489: begin
     mem_space[489] <= din;
    end
    9'd490: begin
     mem_space[490] <= din;
    end
    9'd491: begin
     mem_space[491] <= din;
    end
    9'd492: begin
     mem_space[492] <= din;
    end
    9'd493: begin
     mem_space[493] <= din;
    end
    9'd494: begin
     mem_space[494] <= din;
    end
    9'd495: begin
     mem_space[495] <= din;
    end
    9'd496: begin
     mem_space[496] <= din;
    end
    9'd497: begin
     mem_space[497] <= din;
    end
    9'd498: begin
     mem_space[498] <= din;
    end
    9'd499: begin
     mem_space[499] <= din;
    end
    9'd500: begin
     mem_space[500] <= din;
    end
    9'd501: begin
     mem_space[501] <= din;
    end
    9'd502: begin
     mem_space[502] <= din;
    end
    9'd503: begin
     mem_space[503] <= din;
    end
    9'd504: begin
     mem_space[504] <= din;
    end
    9'd505: begin
     mem_space[505] <= din;
    end
    9'd506: begin
     mem_space[506] <= din;
    end
    9'd507: begin
     mem_space[507] <= din;
    end
    9'd508: begin
     mem_space[508] <= din;
    end
    9'd509: begin
     mem_space[509] <= din;
    end
    9'd510: begin
     mem_space[510] <= din;
    end
    9'd511: begin
     mem_space[511] <= din;
    end
  endcase
end





endmodule
