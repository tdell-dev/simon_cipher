module simon64s96_enc (
  input wire clk,
  input wire rst
  );

  endmodule
