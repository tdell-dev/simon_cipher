//Simon Sim top level
//
module simon_sim_top #(
) (
    
