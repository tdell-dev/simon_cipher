class simon_tester;
