`ifndef SIMON_DEFINES
`define SIMON_DEFINES

  `define ADDER_WIDTH 4
  `define NO_OF_TRANSACTIONS 1000

`endif
