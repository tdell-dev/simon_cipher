module simon48s96_enc (
  input wire clk,
  input wire rst
  );

  endmodule
