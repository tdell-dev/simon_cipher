package simon_pkg;

`include "../src/simon_macros.svh"
`include "./tb_classes/simon_tester.svh"
`include "./tb_classes/simon_scoreboard.svh"
`include "./tb_classes/simon_testbench.svh"

endpackage : simon_pkg
