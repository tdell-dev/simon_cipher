`timescale 1ns / 1ps
package simon_sim_headers;

  `include "simon_cfg_if.sv"

  `include "simon_data_if.sv"

  `include "simon_clk.sv"

endpackage : simon_sim_headers
