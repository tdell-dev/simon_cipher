/home/t/Desktop/xsim_verif_example/Adder_4_bit/src/design/adder_4_bit.sv