`ifndef SIMON_TEST_LIST
`define SIMON_TEST_LIST

package simon_test_list;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import simon_env_pkg::*;
  import simon_seq_list::*;

  //including test list
  `include "simon_basic_test.sv"

endpackage
`endif
