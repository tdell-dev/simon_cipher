module simon64s128_enc (
  input wire clk,
  input wire rst
  );

  endmodule
