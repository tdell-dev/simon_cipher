module simon96s144_enc (
  input wire clk,
  input wire rst
  );

  endmodule
