module simon128s256_enc (
  input wire clk,
  input wire rst
  );

  endmodule
