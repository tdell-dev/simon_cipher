parameter CFG_DATA_WIDTH    =  32;
parameter CFG_ADDR_WIDTH    =  32;
parameter CFG_PROT_WIDTH    =   1;
parameter CFG_RESP_WIDTH    =   2;
parameter CFG_STRB_WIDTH    =   4;

parameter DATA_DATA_WIDTH   = 128;
parameter DATA_ADDR_WIDTH   =  32;
parameter DATA_BURST_WIDTH  =   2;
parameter DATA_CACHE_WIDTH  =   4;
parameter DATA_LEN_WIDTH    =   8;
parameter DATA_LOCK_WIDTH   =   1;
parameter DATA_PROT_WIDTH   =   3;
parameter DATA_QOS_WIDTH    =   4;
parameter DATA_REGION_WIDTH =   4;
parameter DATA_SIZE_WIDTH   =   3;
parameter DATA_RESP_WIDTH   =   2;
parameter DATA_STRB_WIDTH   =  16;
