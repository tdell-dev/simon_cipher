module simon48s72_enc (
  input wire clk,
  input wire rst
  );

  endmodule
